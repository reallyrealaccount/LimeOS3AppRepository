76 69 70 0 0 0 0 0 1 0 0 0 0 0 0 0 57 66 105 116 66 121 116 101 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 50 99 102 99 54 98 101 99 102 54 53 48 49 55 53 52 55 55 57 98 97 50 48 49 99 97 54 52 50 100 97 54 48 49 52 55 53 57 97 48 52 97 56 99 50 57 100 53 101 52 48 57 55 99 99 55 98 98 97 99 49 52 56 49 27 76 117 97 81 0 1 4 8 4 8 0 2 0 0 0 0 0 0 0 64 0 0 0 0 0 0 0 0 0 0 0 2 3 9 0 0 0 5 0 0 0 6 64 64 0 65 128 0 0 28 128 0 1 6 192 64 0 11 0 65 0 164 0 0 0 28 64 128 1 30 0 128 0 5 0 0 0 4 5 0 0 0 0 0 0 0 76 105 109 101 0 4 11 0 0 0 0 0 0 0 71 101 116 83 101 114 118 105 99 101 0 4 11 0 0 0 0 0 0 0 82 117 110 83 101 114 118 105 99 101 0 4 14 0 0 0 0 0 0 0 82 101 110 100 101 114 83 116 101 112 112 101 100 0 4 8 0 0 0 0 0 0 0 67 111 110 110 101 99 116 0 1 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 3 0 0 0 0 0 0 2 5 0 0 0 5 0 0 0 6 64 64 0 65 128 0 0 28 64 0 1 30 0 128 0 3 0 0 0 4 5 0 0 0 0 0 0 0 76 105 109 101 0 4 13 0 0 0 0 0 0 0 67 114 101 97 116 101 87 105 110 100 111 119 0 4 1 0 0 0 0 0 0 0 0 0 0 0 0 5 0 0 0 2 0 0 0 2 0 0 0 2 0 0 0 2 0 0 0 3 0 0 0 0 0 0 0 0 0 0 0 9 0 0 0 1 0 0 0 1 0 0 0 1 0 0 0 1 0 0 0 1 0 0 0 1 0 0 0 3 0 0 0 1 0 0 0 3 0 0 0 0 0 0 0 0 0 0 0 