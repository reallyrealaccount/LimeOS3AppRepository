76 69 70 0 0 0 0 0 1 0 0 0 0 0 0 0 57 66 105 116 66 121 116 101 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 53 54 102 101 100 51 99 101 50 48 50 57 49 51 49 56 97 49 52 54 56 101 55 56 98 52 50 51 55 56 49 97 101 57 56 100 53 57 54 98 102 50 100 98 98 55 49 54 98 52 50 56 99 56 98 55 56 48 57 55 100 100 53 99 27 76 117 97 81 0 1 4 8 4 8 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 2 97 139 5 0 0 5 0 0 0 28 128 128 0 6 64 64 0 69 0 0 0 92 128 128 0 70 128 192 0 133 0 0 0 156 128 128 0 134 192 64 1 197 0 0 0 220 128 128 0 198 0 193 1 0 1 128 0 65 65 1 0 28 129 0 1 70 129 65 0 129 193 1 0 92 129 0 1 134 1 66 2 198 65 66 2 220 129 128 0 1 130 2 0 213 1 130 3 156 129 0 1 154 65 0 0 22 128 1 128 134 193 66 2 198 65 66 2 220 129 128 0 1 130 2 0 213 1 130 3 1 2 3 0 156 65 128 1 134 1 66 2 198 65 66 2 220 129 128 0 1 66 3 0 213 1 130 3 156 129 0 1 154 65 0 0 22 128 1 128 134 193 66 2 198 65 66 2 220 129 128 0 1 66 3 0 213 1 130 3 1 2 3 0 156 65 128 1 134 129 67 0 193 193 3 0 156 129 0 1 195 1 128 3 6 2 68 0 65 66 4 0 128 2 0 3 28 130 128 1 69 194 4 0 70 2 197 4 129 66 5 0 193 66 5 0 92 130 128 1 9 66 2 137 9 194 69 139 70 2 68 0 129 2 6 0 192 2 0 4 92 130 128 1 133 194 4 0 134 2 69 5 193 66 6 0 1 67 6 0 156 130 128 1 73 130 2 137 133 194 4 0 134 2 69 5 193 194 6 0 1 195 6 0 156 130 128 1 73 130 2 141 73 66 71 142 73 194 71 143 73 66 69 144 133 130 8 0 134 194 72 5 193 2 9 0 1 3 9 0 65 3 9 0 156 130 0 2 73 130 130 144 73 130 201 146 134 2 68 0 193 2 6 0 0 3 0 4 156 130 128 1 197 194 4 0 198 2 197 5 1 67 6 0 65 67 6 0 220 130 128 1 137 194 2 137 197 194 4 0 198 2 197 5 1 195 6 0 65 3 9 0 220 130 128 1 137 194 2 141 137 66 71 142 137 194 73 143 137 66 69 144 197 130 8 0 198 194 200 5 1 3 9 0 65 3 9 0 129 3 9 0 220 130 0 2 137 194 130 144 137 130 201 146 198 2 68 0 1 67 4 0 64 3 0 4 220 130 128 1 5 195 4 0 6 3 69 6 65 195 6 0 129 195 6 0 28 131 128 1 201 2 3 137 5 195 4 0 6 3 69 6 65 3 10 0 129 3 10 0 28 131 128 1 201 2 3 141 5 131 8 0 6 195 72 6 65 3 9 0 129 3 9 0 193 3 9 0 28 131 0 2 201 2 131 148 201 194 74 149 201 194 69 139 201 2 203 146 6 3 68 0 65 3 6 0 128 3 128 5 28 131 128 1 69 195 4 0 70 3 197 6 129 195 10 0 193 67 11 0 92 131 128 1 9 67 3 137 69 195 4 0 70 3 197 6 129 131 11 0 193 3 9 0 92 131 128 1 9 67 3 141 9 67 71 142 9 195 75 143 9 67 69 144 69 131 8 0 70 195 200 6 129 3 12 0 193 3 12 0 1 4 12 0 92 131 0 2 9 67 131 144 70 3 68 0 129 67 12 0 192 3 128 5 92 131 128 1 133 195 4 0 134 3 69 7 193 131 12 0 1 132 11 0 156 131 128 1 73 131 3 137 133 195 4 0 134 3 69 7 193 67 6 0 1 68 11 0 156 131 128 1 73 131 3 141 73 67 71 142 73 195 76 143 73 3 77 144 133 131 8 0 134 195 72 7 193 3 12 0 1 4 12 0 65 4 12 0 156 131 0 2 73 131 131 144 134 3 68 0 193 67 12 0 0 4 128 5 156 131 128 1 197 195 4 0 198 3 197 7 1 68 13 0 65 132 11 0 220 131 128 1 137 195 3 137 197 195 4 0 198 3 197 7 1 68 6 0 65 132 13 0 220 131 128 1 137 195 3 141 137 67 71 142 137 195 77 143 137 3 77 144 197 131 8 0 198 195 200 7 1 4 12 0 65 4 12 0 129 4 12 0 220 131 0 2 137 195 131 144 198 3 68 0 1 68 12 0 64 4 128 5 220 131 128 1 5 196 4 0 6 4 69 8 65 68 13 0 129 132 11 0 28 132 128 1 201 3 4 137 5 196 4 0 6 4 69 8 65 4 14 0 129 132 13 0 28 132 128 1 201 3 4 141 201 67 71 142 201 67 78 143 201 3 77 144 5 132 8 0 6 196 72 8 65 4 12 0 129 4 12 0 193 4 12 0 28 132 0 2 201 3 132 144 6 4 68 0 65 68 12 0 128 4 128 5 28 132 128 1 69 196 4 0 70 4 197 8 129 132 12 0 193 132 11 0 92 132 128 1 9 68 4 137 69 196 4 0 70 4 197 8 129 68 6 0 193 132 14 0 92 132 128 1 9 68 4 141 9 68 71 142 9 196 78 143 9 4 77 144 69 132 8 0 70 196 200 8 129 4 12 0 193 4 12 0 1 5 12 0 92 132 0 2 9 68 132 144 70 4 68 0 129 68 4 0 192 4 0 3 92 132 128 1 133 196 4 0 134 4 69 9 193 68 5 0 1 69 5 0 156 132 128 1 73 132 4 137 134 4 68 0 193 68 4 0 0 5 0 3 156 132 128 1 197 196 4 0 198 4 197 9 1 69 5 0 65 69 5 0 220 132 128 1 137 196 4 137 137 196 69 139 198 4 68 0 1 5 15 0 64 5 0 9 220 132 128 1 201 68 79 143 201 196 79 159 5 197 4 0 6 5 69 10 65 197 10 0 129 133 11 0 28 133 128 1 201 4 5 137 5 197 4 0 6 5 69 10 65 133 11 0 129 5 10 0 28 133 128 1 201 4 5 141 6 5 68 0 65 69 4 0 128 5 0 3 28 133 128 1 69 197 4 0 70 5 197 10 129 69 5 0 193 69 5 0 92 133 128 1 9 69 5 137 9 197 69 139 70 5 68 0 129 5 16 0 192 5 0 10 92 133 128 1 133 197 4 0 134 5 69 11 193 197 6 0 1 70 16 0 156 133 128 1 73 133 5 137 133 197 4 0 134 5 69 11 193 5 10 0 1 6 9 0 156 133 128 1 73 133 5 141 133 197 16 0 134 5 81 11 134 69 81 11 73 133 5 161 134 5 68 0 193 133 17 0 0 6 128 10 156 69 128 1 134 5 68 0 193 69 12 0 0 6 0 10 156 133 128 1 197 197 4 0 198 5 197 11 1 70 13 0 65 198 17 0 220 133 128 1 137 197 5 137 197 197 4 0 198 5 197 11 1 6 10 0 65 6 18 0 220 133 128 1 137 197 5 141 137 69 71 142 137 69 82 143 137 5 77 144 197 133 8 0 198 197 200 11 1 6 12 0 65 6 12 0 129 6 12 0 220 133 0 2 137 197 133 144 198 5 68 0 1 70 12 0 64 6 0 10 220 133 128 1 5 198 4 0 6 6 69 12 65 70 13 0 129 198 17 0 28 134 128 1 201 5 6 137 5 198 4 0 6 6 69 12 65 6 14 0 129 6 18 0 28 134 128 1 201 5 6 141 201 69 71 142 201 133 82 143 201 5 77 144 5 134 8 0 6 198 72 12 65 6 12 0 129 6 12 0 193 6 12 0 28 134 0 2 201 5 134 144 6 6 68 0 65 70 4 0 128 6 0 3 28 134 128 1 69 198 4 0 70 6 197 12 129 70 5 0 193 70 5 0 92 134 128 1 9 70 6 137 9 198 69 139 70 6 68 0 129 70 4 0 192 6 0 3 92 134 128 1 133 198 4 0 134 6 69 13 193 70 5 0 1 71 5 0 156 134 128 1 73 134 6 137 73 198 69 139 134 6 68 0 193 6 6 0 0 7 128 12 156 134 128 1 197 198 4 0 198 6 197 13 1 199 10 0 65 71 11 0 220 134 128 1 137 198 6 137 197 198 4 0 198 6 197 13 1 135 11 0 65 7 9 0 220 134 128 1 137 198 6 141 137 70 71 142 137 198 82 143 137 70 69 144 197 134 8 0 198 198 200 13 1 7 12 0 65 7 12 0 129 7 12 0 220 134 0 2 137 198 134 144 198 6 68 0 1 7 15 0 64 7 0 12 220 134 128 1 5 199 4 0 6 7 69 14 65 71 13 0 129 135 11 0 28 135 128 1 201 6 7 137 5 199 4 0 6 7 69 14 65 7 10 0 129 7 9 0 28 135 128 1 201 6 7 141 201 70 71 142 201 6 83 143 201 70 83 159 201 198 74 144 5 135 8 0 6 199 72 14 65 7 12 0 129 7 12 0 193 7 12 0 28 135 0 2 201 6 135 144 6 7 68 0 65 7 15 0 128 7 0 12 28 135 128 1 69 199 4 0 70 7 197 14 129 71 13 0 193 135 11 0 92 135 128 1 9 71 7 137 69 199 4 0 70 7 197 14 129 7 14 0 193 7 9 0 92 135 128 1 9 71 7 141 9 71 71 142 9 7 83 143 9 135 83 159 9 199 74 144 69 135 8 0 70 199 200 14 129 7 12 0 193 7 12 0 1 8 12 0 92 135 0 2 9 71 135 144 70 7 68 0 129 7 15 0 192 7 0 12 92 135 128 1 133 199 4 0 134 7 69 15 193 71 11 0 1 136 11 0 156 135 128 1 73 135 7 137 133 199 4 0 134 7 69 15 193 7 10 0 1 200 19 0 156 135 128 1 73 135 7 141 73 71 71 142 73 7 84 143 73 71 84 159 73 199 74 144 133 135 8 0 134 199 72 15 193 7 12 0 1 8 12 0 65 8 12 0 156 135 0 2 73 135 135 144 134 7 68 0 193 7 15 0 0 8 0 12 156 135 128 1 197 199 4 0 198 7 197 15 1 72 11 0 65 136 11 0 220 135 128 1 137 199 7 137 197 199 4 0 198 7 197 15 1 136 20 0 65 200 19 0 220 135 128 1 137 199 7 141 137 71 71 142 137 7 84 143 137 199 84 159 137 199 74 144 197 135 8 0 198 199 200 15 1 8 12 0 65 8 12 0 129 8 12 0 220 135 0 2 137 199 135 144 198 7 68 0 1 8 15 0 64 8 0 12 220 135 128 1 5 200 4 0 6 8 69 16 65 72 11 0 129 136 11 0 28 136 128 1 201 7 8 137 5 200 4 0 6 8 69 16 65 8 21 0 129 200 19 0 28 136 128 1 201 7 8 141 201 71 71 142 201 71 85 143 201 135 85 159 201 199 74 144 5 136 8 0 6 200 72 16 65 8 12 0 129 8 12 0 193 8 12 0 28 136 0 2 201 7 136 144 6 8 68 0 65 72 12 0 128 8 0 12 28 136 128 1 69 200 4 0 70 8 197 16 129 200 10 0 193 136 11 0 92 136 128 1 9 72 8 137 69 200 4 0 70 8 197 16 129 136 11 0 193 200 10 0 92 136 128 1 9 72 8 141 9 72 71 142 9 200 85 143 9 200 74 144 69 136 8 0 70 200 200 16 129 8 12 0 193 8 12 0 1 9 12 0 92 136 0 2 9 72 136 144 70 8 68 0 129 72 12 0 192 8 0 9 92 136 128 1 133 200 4 0 134 8 69 17 193 72 13 0 1 137 11 0 156 136 128 1 73 136 8 137 133 200 4 0 134 8 69 17 193 72 11 0 1 137 14 0 156 136 128 1 73 136 8 141 73 72 71 142 73 8 86 143 73 8 77 144 133 136 8 0 134 200 72 17 193 8 12 0 1 9 12 0 65 9 12 0 156 136 0 2 73 136 136 144 134 8 68 0 193 72 22 0 0 9 128 8 156 136 128 1 197 200 4 0 198 8 197 17 1 73 5 0 65 73 5 0 220 136 128 1 137 200 8 137 137 72 69 144 198 8 68 0 1 9 6 0 64 9 128 8 220 136 128 1 5 201 4 0 6 9 69 18 65 73 16 0 129 73 11 0 28 137 128 1 201 8 9 137 5 201 4 0 6 9 69 18 65 73 6 0 129 9 9 0 28 137 128 1 201 8 9 141 201 72 71 142 201 200 67 143 201 72 69 144 5 137 8 0 6 201 72 18 65 9 12 0 129 9 12 0 193 9 12 0 28 137 0 2 201 8 137 144 6 9 68 0 65 73 12 0 128 9 128 8 28 137 128 1 69 201 4 0 70 9 197 18 129 73 16 0 193 137 11 0 92 137 128 1 9 73 9 137 69 201 4 0 70 9 197 18 129 73 6 0 193 73 11 0 92 137 128 1 9 73 9 141 9 73 71 142 9 137 86 143 9 9 77 144 69 137 8 0 70 201 200 18 129 9 12 0 193 9 12 0 1 10 12 0 92 137 0 2 9 73 137 144 70 9 68 0 129 73 12 0 192 9 128 8 92 137 128 1 133 201 4 0 134 9 69 19 193 73 13 0 1 138 11 0 156 137 128 1 73 137 9 137 133 201 4 0 134 9 69 19 193 73 6 0 1 138 13 0 156 137 128 1 73 137 9 141 73 73 71 142 73 73 78 143 73 9 77 144 133 137 8 0 134 201 72 19 193 9 12 0 1 10 12 0 65 10 12 0 156 137 0 2 73 137 137 144 134 9 68 0 193 73 12 0 0 10 128 8 156 137 128 1 197 201 4 0 198 9 197 19 1 74 13 0 65 138 11 0 220 137 128 1 137 201 9 137 197 201 4 0 198 9 197 19 1 202 22 0 65 138 13 0 220 137 128 1 137 201 9 141 137 73 71 142 137 9 87 143 137 9 77 144 197 137 8 0 198 201 200 19 1 10 12 0 65 10 12 0 129 10 12 0 220 137 0 2 137 201 137 144 198 9 68 0 1 74 12 0 64 10 128 8 220 137 128 1 5 202 4 0 6 10 69 20 65 74 16 0 129 138 11 0 28 138 128 1 201 9 10 137 5 202 4 0 6 10 69 20 65 74 6 0 129 138 14 0 28 138 128 1 201 9 10 141 201 73 71 142 201 73 87 143 201 9 77 144 5 138 8 0 6 202 72 20 65 10 12 0 129 10 12 0 193 10 12 0 28 138 0 2 201 9 138 144 6 10 68 0 65 74 4 0 128 10 0 3 28 138 128 1 69 202 4 0 70 10 197 20 129 74 5 0 193 74 5 0 92 138 128 1 9 74 10 137 9 202 69 139 70 10 68 0 129 10 6 0 192 10 0 20 92 138 128 1 133 202 4 0 134 10 69 21 193 74 5 0 1 75 16 0 156 138 128 1 73 138 10 137 73 74 71 142 73 10 77 144 73 138 87 143 133 138 8 0 134 202 72 21 193 10 12 0 1 11 12 0 65 11 12 0 156 138 0 2 73 138 138 144 134 10 68 0 193 74 12 0 0 11 0 20 156 138 128 1 197 202 4 0 198 10 197 21 1 75 5 0 65 139 11 0 220 138 128 1 137 202 10 137 197 202 4 0 198 10 197 21 1 11 9 0 65 75 16 0 220 138 128 1 137 202 10 141 137 74 71 142 137 10 77 144 137 10 86 143 197 138 8 0 198 202 200 21 1 11 12 0 65 11 12 0 129 11 12 0 220 138 0 2 137 202 138 144 198 202 215 19 203 10 216 21 100 11 0 0 0 0 128 0 0 0 0 3 220 74 128 1 198 202 215 18 203 10 216 21 100 75 0 0 0 0 128 8 0 0 0 4 0 0 128 12 0 0 0 9 220 74 128 1 198 202 87 19 203 10 216 21 100 139 0 0 0 0 128 8 0 0 0 4 0 0 128 12 0 0 0 20 220 74 128 1 198 202 87 21 203 10 216 21 100 203 0 0 0 0 0 20 0 0 0 9 0 0 128 5 0 0 128 8 0 0 0 4 220 74 128 1 198 202 215 16 203 10 216 21 100 11 1 0 0 0 128 12 0 0 0 9 0 0 128 5 0 0 128 8 0 0 0 4 220 74 128 1 198 202 215 7 203 10 216 21 100 75 1 0 0 0 128 8 0 0 0 4 0 0 128 12 0 0 0 9 220 74 128 1 198 10 68 0 1 75 24 0 64 11 0 4 220 138 128 1 5 203 4 0 6 11 69 22 65 75 5 0 129 75 5 0 28 139 128 1 201 10 11 137 5 139 8 0 6 203 72 22 65 75 15 0 129 75 15 0 193 75 15 0 28 139 0 2 201 10 11 177 6 203 216 9 11 11 88 22 164 139 1 0 0 0 128 21 0 0 128 9 28 75 128 1 6 11 68 0 65 11 25 0 128 11 128 21 28 139 128 1 70 11 68 0 129 75 25 0 192 11 0 22 92 139 128 1 134 11 68 0 193 11 6 0 0 12 0 4 156 139 128 1 197 203 4 0 198 11 197 23 1 76 6 0 65 76 6 0 220 139 128 1 137 203 11 137 137 139 89 143 137 75 71 142 197 139 8 0 198 203 200 23 1 12 12 0 65 12 12 0 129 12 12 0 220 139 0 2 137 203 139 144 137 75 69 144 197 203 4 0 198 11 197 23 1 204 25 0 65 204 25 0 220 139 128 1 137 203 11 141 198 11 68 0 1 12 6 0 64 12 0 4 220 139 128 1 5 204 4 0 6 12 69 24 65 76 6 0 129 76 6 0 28 140 128 1 201 11 12 137 201 75 71 142 201 75 69 144 5 140 8 0 6 204 72 24 65 12 9 0 129 12 9 0 193 12 9 0 28 140 0 2 201 11 140 144 201 11 90 143 1 76 26 0 65 76 26 0 129 140 26 0 193 204 26 0 1 13 27 0 100 205 1 0 0 0 0 24 0 0 0 25 0 0 128 24 0 0 0 0 0 0 128 22 164 13 2 0 0 0 0 25 0 0 128 25 0 0 0 26 0 0 128 26 193 13 11 0 1 78 27 0 74 14 128 4 138 142 0 0 197 206 27 0 198 14 220 29 1 15 9 0 65 79 5 0 129 15 9 0 220 142 0 2 137 206 14 183 197 142 8 0 198 206 200 29 1 143 28 0 65 207 28 0 129 15 29 0 220 142 0 2 137 206 142 184 202 142 0 0 5 207 27 0 6 15 92 30 65 15 9 0 129 143 26 0 193 15 9 0 28 143 0 2 201 14 15 183 5 143 8 0 6 207 72 30 65 143 28 0 129 207 28 0 193 15 29 0 28 143 0 2 201 14 143 184 10 143 0 0 69 207 27 0 70 15 220 30 129 15 9 0 193 79 29 0 1 16 9 0 92 143 0 2 9 79 15 183 69 143 8 0 70 207 200 30 129 143 28 0 193 207 28 0 1 16 29 0 92 143 0 2 9 79 143 184 74 143 0 0 133 207 27 0 134 15 92 31 193 15 9 0 1 144 29 0 65 16 9 0 156 143 0 2 73 143 15 183 133 143 8 0 134 207 72 31 193 143 28 0 1 208 28 0 65 16 29 0 156 143 0 2 73 143 143 184 138 143 0 0 197 207 27 0 198 15 220 31 1 16 9 0 65 208 29 0 129 16 9 0 220 143 0 2 137 207 15 183 197 143 8 0 198 207 200 31 1 16 30 0 65 80 30 0 129 16 9 0 220 143 0 2 137 207 143 184 202 143 0 0 5 208 27 0 6 16 92 32 65 80 5 0 129 144 29 0 193 16 9 0 28 144 0 2 201 15 16 183 5 144 8 0 6 208 72 32 65 16 30 0 129 80 30 0 193 16 9 0 28 144 0 2 201 15 144 184 10 144 0 0 69 208 27 0 70 16 220 32 129 144 30 0 193 144 29 0 1 17 9 0 92 144 0 2 9 80 16 183 69 144 8 0 70 208 200 32 129 16 30 0 193 80 30 0 1 17 9 0 92 144 0 2 9 80 144 184 74 144 0 0 133 208 27 0 134 16 92 33 193 16 9 0 1 145 29 0 65 81 5 0 156 144 0 2 73 144 16 183 133 144 8 0 134 208 72 33 193 16 30 0 1 81 30 0 65 17 9 0 156 144 0 2 73 144 144 184 138 144 0 0 197 208 27 0 198 16 220 33 1 17 9 0 65 145 29 0 129 145 30 0 220 144 0 2 137 208 16 183 197 144 8 0 198 208 200 33 1 17 30 0 65 81 30 0 129 17 9 0 220 144 0 2 137 208 144 184 98 78 128 4 138 14 0 0 228 78 2 0 0 0 128 24 0 0 0 24 0 0 128 27 0 0 0 27 0 0 0 28 0 0 0 25 0 0 128 25 0 0 0 26 0 0 128 28 0 0 0 29 0 0 128 26 0 0 0 13 6 15 68 0 65 207 30 0 128 15 0 22 28 143 128 1 201 10 15 190 9 143 223 190 65 15 9 0 129 15 9 0 193 207 31 0 6 144 65 0 65 16 32 0 28 144 0 1 64 16 128 1 92 144 128 0 164 144 2 0 0 0 0 32 0 0 128 30 0 0 128 31 0 0 0 31 0 0 0 30 135 80 32 0 138 16 0 3 197 144 8 0 198 208 200 33 1 17 30 0 65 81 30 0 129 17 9 0 220 144 0 2 5 145 8 0 6 209 72 34 65 145 28 0 129 209 28 0 193 17 29 0 28 145 0 2 69 145 8 0 70 209 200 34 129 145 32 0 193 145 32 0 1 146 32 0 92 145 0 2 133 145 8 0 134 209 72 35 193 17 9 0 1 18 9 0 65 210 32 0 156 145 0 2 197 145 8 0 198 209 200 35 1 18 9 0 65 18 33 0 129 82 33 0 220 145 0 2 5 146 8 0 6 210 72 36 65 146 33 0 129 210 33 0 193 18 34 0 28 146 0 2 69 146 8 0 70 210 200 36 129 18 12 0 193 18 12 0 1 19 12 0 92 18 0 2 162 80 0 0 193 80 34 0 36 209 2 0 0 0 0 25 0 0 128 33 0 0 0 1 100 17 3 0 0 0 0 1 0 0 128 26 0 0 0 25 0 0 128 33 0 0 0 24 71 145 34 0 100 81 3 0 0 0 0 33 0 0 0 24 0 0 128 24 0 0 128 33 164 145 3 0 0 0 0 24 0 0 128 24 0 0 128 33 0 0 0 33 228 209 3 0 0 0 0 2 0 0 128 22 0 0 128 34 0 0 0 34 36 18 4 0 0 0 0 2 0 0 0 35 78 146 140 187 134 18 68 0 193 82 12 0 0 19 0 4 156 146 128 1 137 210 226 146 137 82 69 144 137 18 83 143 197 210 4 0 198 18 197 37 1 83 5 0 65 83 5 0 220 146 128 1 137 210 18 137 195 18 128 38 164 83 4 0 0 0 0 22 0 0 0 30 0 0 128 36 228 147 4 0 0 0 0 22 0 0 0 30 0 0 128 36 0 0 0 25 0 0 128 26 6 20 99 37 11 20 88 40 164 212 4 0 0 0 0 32 0 0 0 39 28 84 128 1 6 84 99 37 11 20 88 40 164 20 5 0 0 0 0 32 0 0 128 39 28 84 128 1 6 148 227 32 11 20 88 40 164 84 5 0 0 0 0 32 0 0 0 39 28 148 128 1 0 19 0 40 6 212 227 32 11 20 88 40 164 148 5 0 0 0 0 32 0 0 128 39 28 148 128 1 64 19 0 40 36 212 5 0 0 0 0 0 0 0 128 2 70 20 100 32 75 20 216 40 228 20 6 0 0 0 0 4 0 0 0 32 0 0 128 5 0 0 0 37 0 0 0 30 0 0 0 40 92 148 128 1 192 18 128 40 70 212 215 6 75 20 216 40 228 84 6 0 0 0 0 32 0 0 0 37 0 0 128 5 92 84 128 1 70 212 87 8 75 20 216 40 228 148 6 0 0 0 128 22 0 0 0 0 0 0 0 22 0 0 128 3 0 0 0 4 0 0 128 5 0 0 128 8 92 84 128 1 70 84 228 32 75 20 216 40 197 84 32 0 92 84 128 1 65 148 36 0 129 212 22 0 193 20 9 0 14 149 140 201 18 21 0 42 65 149 12 0 142 149 12 202 206 149 140 202 36 214 6 0 0 0 0 22 100 22 7 0 0 0 0 44 0 0 0 30 0 0 0 41 164 86 7 0 0 0 0 0 0 0 128 3 0 0 0 32 0 0 0 30 0 0 128 44 0 0 0 43 0 0 0 22 0 0 128 40 0 0 128 43 0 0 128 41 0 0 0 25 0 0 0 42 0 0 128 42 0 0 128 23 0 0 0 5 193 22 19 0 6 215 87 18 11 23 88 46 164 151 7 0 0 0 128 8 0 0 0 4 0 0 128 12 0 0 0 9 0 0 0 10 0 0 128 10 0 0 0 2 0 0 0 0 0 0 128 45 28 87 128 1 36 215 7 0 0 0 0 32 0 0 0 1 0 0 0 4 0 0 128 12 0 0 0 10 0 0 0 12 0 0 0 45 0 0 0 30 0 0 0 25 65 23 19 0 134 215 215 11 139 23 88 47 36 24 8 0 0 0 128 45 0 0 128 46 0 0 0 36 0 0 0 46 156 87 128 1 134 215 87 11 139 23 88 47 36 88 8 0 0 0 0 10 0 0 0 12 156 87 128 1 134 215 87 16 139 23 88 47 36 152 8 0 0 0 0 12 0 0 128 12 0 0 128 46 0 0 0 14 0 0 0 24 0 0 128 14 0 0 128 24 0 0 0 15 0 0 128 15 0 0 128 33 0 0 0 25 0 0 128 29 0 0 128 13 0 0 0 46 156 87 128 1 134 215 87 7 139 23 88 47 36 216 8 0 0 0 128 35 0 0 128 46 0 0 0 32 0 0 0 37 0 0 128 5 156 87 128 1 128 23 128 0 193 151 37 0 156 151 0 1 134 215 101 47 198 23 102 3 198 87 230 47 198 87 230 47 36 24 9 0 0 0 0 1 0 0 128 3 0 0 128 37 0 0 0 38 0 0 128 38 156 87 128 1 30 0 128 0 154 0 0 0 4 8 0 0 0 0 0 0 0 103 101 116 102 101 110 118 0 4 5 0 0 0 0 0 0 0 76 105 109 101 0 4 8 0 0 0 0 0 0 0 108 111 97 100 108 105 98 0 4 4 0 0 0 0 0 0 0 108 111 103 0 4 9 0 0 0 0 0 0 0 71 101 116 77 111 117 115 101 0 4 11 0 0 0 0 0 0 0 70 105 108 101 83 121 115 116 101 109 0 4 11 0 0 0 0 0 0 0 71 101 116 83 101 114 118 105 99 101 0 4 13 0 0 0 0 0 0 0 83 111 117 110 100 83 101 114 118 105 99 101 0 4 11 0 0 0 0 0 0 0 70 105 108 101 69 120 105 115 116 115 0 4 17 0 0 0 0 0 0 0 71 101 116 79 83 68 114 105 118 101 76 101 116 116 101 114 0 4 28 0 0 0 0 0 0 0 58 47 83 121 115 116 101 109 47 65 112 112 68 97 116 97 47 66 117 105 108 100 66 114 101 97 107 0 4 16 0 0 0 0 0 0 0 67 114 101 97 116 101 68 105 114 101 99 116 111 114 121 0 4 8 0 0 0 0 0 0 0 82 45 87 45 68 45 65 0 4 34 0 0 0 0 0 0 0 58 47 83 121 115 116 101 109 47 65 112 112 68 97 116 97 47 66 117 105 108 100 66 114 101 97 107 47 115 97 118 101 115 0 4 13 0 0 0 0 0 0 0 67 114 101 97 116 101 87 105 110 100 111 119 0 4 11 0 0 0 0 0 0 0 66 117 105 108 100 66 114 101 97 107 0 4 9 0 0 0 0 0 0 0 67 114 101 97 116 101 85 73 0 4 6 0 0 0 0 0 0 0 70 114 97 109 101 0 4 5 0 0 0 0 0 0 0 83 105 122 101 0 4 6 0 0 0 0 0 0 0 85 68 105 109 50 0 4 10 0 0 0 0 0 0 0 102 114 111 109 83 99 97 108 101 0 3 0 0 0 0 0 0 240 63 4 8 0 0 0 0 0 0 0 86 105 115 105 98 108 101 0 1 0 4 10 0 0 0 0 0 0 0 84 101 120 116 76 97 98 101 108 0 3 154 153 153 153 153 153 185 63 4 9 0 0 0 0 0 0 0 80 111 115 105 116 105 111 110 0 3 205 204 204 204 204 204 236 63 4 11 0 0 0 0 0 0 0 84 101 120 116 83 99 97 108 101 100 0 1 1 4 5 0 0 0 0 0 0 0 84 101 120 116 0 4 15 0 0 0 0 0 0 0 118 48 46 50 46 48 32 114 101 108 101 97 115 101 0 4 23 0 0 0 0 0 0 0 66 97 99 107 103 114 111 117 110 100 84 114 97 110 115 112 97 114 101 110 99 121 0 4 11 0 0 0 0 0 0 0 84 101 120 116 67 111 108 111 114 51 0 4 7 0 0 0 0 0 0 0 67 111 108 111 114 51 0 4 8 0 0 0 0 0 0 0 102 114 111 109 82 71 66 0 3 0 0 0 0 0 0 0 0 4 7 0 0 0 0 0 0 0 90 73 110 100 101 120 0 3 0 0 0 0 0 0 38 64 4 6 0 0 0 0 0 0 0 88 32 89 32 90 0 3 154 153 153 153 153 153 169 63 4 17 0 0 0 0 0 0 0 66 97 99 107 103 114 111 117 110 100 67 111 108 111 114 51 0 4 13 0 0 0 0 0 0 0 84 114 97 110 115 112 97 114 101 110 99 121 0 3 51 51 51 51 51 51 227 63 3 0 0 0 0 0 0 36 64 3 51 51 51 51 51 51 211 63 3 154 153 153 153 153 153 201 63 4 7 0 0 0 0 0 0 0 80 97 117 115 101 100 0 3 0 0 0 0 0 224 111 64 4 11 0 0 0 0 0 0 0 84 101 120 116 66 117 116 116 111 110 0 3 51 51 51 51 51 51 235 63 4 13 0 0 0 0 0 0 0 66 97 99 107 32 116 111 32 103 97 109 101 0 3 102 102 102 102 102 102 230 63 3 154 153 153 153 153 153 217 63 3 205 204 204 204 204 204 224 63 4 5 0 0 0 0 0 0 0 83 97 118 101 0 3 154 153 153 153 153 153 225 63 4 9 0 0 0 0 0 0 0 83 101 116 116 105 110 103 115 0 3 0 0 0 0 0 0 232 63 4 15 0 0 0 0 0 0 0 82 101 116 117 114 110 32 116 111 32 109 101 110 117 0 4 8 0 0 0 0 0 0 0 84 101 120 116 66 111 120 0 3 0 0 0 0 0 0 89 64 4 16 0 0 0 0 0 0 0 80 108 97 99 101 104 111 108 100 101 114 84 101 120 116 0 4 6 0 0 0 0 0 0 0 48 45 50 53 53 0 4 15 0 0 0 0 0 0 0 83 99 114 111 108 108 105 110 103 70 114 97 109 101 0 3 154 153 153 153 153 153 233 63 4 20 0 0 0 0 0 0 0 65 117 116 111 109 97 116 105 99 67 97 110 118 97 115 83 105 122 101 0 4 5 0 0 0 0 0 0 0 69 110 117 109 0 4 14 0 0 0 0 0 0 0 65 117 116 111 109 97 116 105 99 83 105 122 101 0 4 2 0 0 0 0 0 0 0 89 0 4 13 0 0 0 0 0 0 0 85 73 76 105 115 116 76 97 121 111 117 116 0 3 51 51 51 51 51 51 195 63 3 102 102 102 102 102 102 234 63 4 9 0 0 0 0 0 0 0 78 101 119 32 103 97 109 101 0 4 10 0 0 0 0 0 0 0 76 111 97 100 32 103 97 109 101 0 4 11 0 0 0 0 0 0 0 76 111 97 100 105 110 103 46 46 46 0 4 1 0 0 0 0 0 0 0 0 4 5 0 0 0 0 0 0 0 83 101 101 100 0 4 10 0 0 0 0 0 0 0 83 97 118 101 32 110 97 109 101 0 3 0 0 0 0 0 0 208 63 4 3 0 0 0 0 0 0 0 52 53 0 4 12 0 0 0 0 0 0 0 87 111 114 108 100 32 119 105 100 116 104 0 3 102 102 102 102 102 102 214 63 4 12 0 0 0 0 0 0 0 87 111 114 108 100 32 100 101 112 116 104 0 3 205 204 204 204 204 204 228 63 4 3 0 0 0 0 0 0 0 54 48 0 4 17 0 0 0 0 0 0 0 87 111 114 108 100 32 109 97 120 32 104 101 105 103 104 116 0 4 5 0 0 0 0 0 0 0 80 108 97 121 0 4 5 0 0 0 0 0 0 0 66 97 99 107 0 4 11 0 0 0 0 0 0 0 73 109 97 103 101 76 97 98 101 108 0 4 6 0 0 0 0 0 0 0 80 108 97 121 33 0 3 0 0 0 0 0 0 224 63 4 9 0 0 0 0 0 0 0 67 111 110 116 114 111 108 115 0 4 5 0 0 0 0 0 0 0 81 117 105 116 0 4 84 0 0 0 0 0 0 0 84 97 98 32 102 111 114 32 112 97 117 115 101 44 32 87 65 83 68 32 116 111 32 109 111 118 101 44 32 109 111 117 115 101 32 116 111 32 108 111 111 107 32 97 114 111 117 110 100 44 32 82 32 116 111 32 114 101 115 101 116 32 112 111 115 105 116 105 111 110 44 32 69 32 102 111 114 32 115 116 101 118 101 0 4 18 0 0 0 0 0 0 0 77 111 117 115 101 66 117 116 116 111 110 49 67 108 105 99 107 0 4 8 0 0 0 0 0 0 0 67 111 110 110 101 99 116 0 4 14 0 0 0 0 0 0 0 86 105 101 119 112 111 114 116 70 114 97 109 101 0 4 8 0 0 0 0 0 0 0 65 109 98 105 101 110 116 0 4 10 0 0 0 0 0 0 0 70 111 99 117 115 76 111 115 116 0 4 11 0 0 0 0 0 0 0 87 111 114 108 100 77 111 100 101 108 0 4 7 0 0 0 0 0 0 0 70 111 108 100 101 114 0 4 2 0 0 0 0 0 0 0 43 0 3 205 204 204 204 204 204 220 63 4 4 0 0 0 0 0 0 0 70 80 83 0 3 0 0 0 0 0 128 70 64 3 0 0 0 0 0 0 0 64 3 0 0 0 0 0 0 78 64 3 0 0 0 0 0 0 68 64 3 0 0 0 0 0 0 105 64 4 4 0 0 0 0 0 0 0 80 111 115 0 4 8 0 0 0 0 0 0 0 86 101 99 116 111 114 51 0 4 4 0 0 0 0 0 0 0 110 101 119 0 4 6 0 0 0 0 0 0 0 67 111 108 111 114 0 3 0 0 0 0 0 0 107 64 3 0 0 0 0 0 160 102 64 3 0 0 0 0 0 32 97 64 3 0 0 0 0 0 0 8 64 3 0 0 0 0 0 0 16 64 3 0 0 0 0 0 0 20 64 3 0 0 0 0 0 0 72 64 3 0 0 0 0 0 224 102 64 3 0 0 0 0 0 0 240 191 4 7 0 0 0 0 0 0 0 67 97 109 101 114 97 0 4 14 0 0 0 0 0 0 0 67 117 114 114 101 110 116 67 97 109 101 114 97 0 4 11 0 0 0 0 0 0 0 67 97 109 101 114 97 84 121 112 101 0 4 11 0 0 0 0 0 0 0 83 99 114 105 112 116 97 98 108 101 0 3 0 0 0 0 0 0 224 191 4 17 0 0 0 0 0 0 0 85 115 101 114 73 110 112 117 116 83 101 114 118 105 99 101 0 4 10 0 0 0 0 0 0 0 77 111 117 115 101 77 111 118 101 0 3 0 0 0 0 0 0 62 64 3 0 0 0 0 0 192 98 64 3 0 0 0 0 0 64 99 64 3 0 0 0 0 0 0 55 64 3 0 0 0 0 0 128 100 64 3 0 0 0 0 0 0 93 64 3 0 0 0 0 0 64 82 64 3 0 0 0 0 0 0 94 64 4 11 0 0 0 0 0 0 0 86 82 76 69 100 101 99 111 100 101 0 3 0 0 0 0 0 56 143 64 4 17 0 0 0 0 0 0 0 77 111 117 115 101 66 117 116 116 111 110 49 68 111 119 110 0 4 17 0 0 0 0 0 0 0 77 111 117 115 101 66 117 116 116 111 110 50 68 111 119 110 0 4 12 0 0 0 0 0 0 0 66 117 116 116 111 110 49 68 111 119 110 0 4 12 0 0 0 0 0 0 0 66 117 116 116 111 110 50 68 111 119 110 0 4 11 0 0 0 0 0 0 0 73 110 112 117 116 66 101 103 97 110 0 4 5 0 0 0 0 0 0 0 77 111 118 101 0 3 123 20 174 71 225 122 132 63 3 154 153 153 153 153 153 35 64 3 248 83 227 165 155 68 17 64 3 0 0 0 0 0 0 248 63 4 19 0 0 0 0 0 0 0 65 112 112 108 105 99 97 116 105 111 110 72 97 110 100 108 101 114 0 4 7 0 0 0 0 0 0 0 79 110 69 120 105 116 0 4 7 0 0 0 0 0 0 0 80 97 114 101 110 116 0 4 6 0 0 0 0 0 0 0 86 97 108 117 101 0 37 0 0 0 0 0 0 0 0 0 0 0 15 1 0 0 17 1 0 0 2 0 0 2 9 0 0 0 4 0 0 0 65 0 0 0 28 128 0 1 6 64 64 0 6 128 64 0 68 0 128 0 70 192 192 0 28 64 0 1 30 0 128 0 4 0 0 0 4 19 0 0 0 0 0 0 0 65 112 112 108 105 99 97 116 105 111 110 72 97 110 100 108 101 114 0 4 5 0 0 0 0 0 0 0 85 115 101 114 0 4 10 0 0 0 0 0 0 0 67 108 111 115 101 80 114 111 99 0 4 7 0 0 0 0 0 0 0 80 97 114 101 110 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 19 1 0 0 24 1 0 0 4 0 0 2 9 0 0 0 4 0 0 0 9 64 64 128 4 0 128 0 9 64 64 128 4 0 0 1 9 64 64 128 4 0 128 1 9 128 64 128 30 0 128 0 3 0 0 0 4 8 0 0 0 0 0 0 0 86 105 115 105 98 108 101 0 1 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 26 1 0 0 31 1 0 0 4 0 0 2 9 0 0 0 4 0 0 0 9 64 64 128 4 0 128 0 9 64 64 128 4 0 0 1 9 64 64 128 4 0 128 1 9 128 64 128 30 0 128 0 3 0 0 0 4 8 0 0 0 0 0 0 0 86 105 115 105 98 108 101 0 1 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 33 1 0 0 43 1 0 0 5 0 0 2 18 0 0 0 4 0 0 0 9 64 64 128 4 0 128 0 9 64 64 128 4 0 0 1 6 0 64 0 26 0 0 0 22 0 1 128 4 0 128 1 9 64 64 128 4 0 0 2 9 128 64 128 22 192 0 128 4 0 128 1 9 128 64 128 4 0 0 2 9 64 64 128 30 0 128 0 3 0 0 0 4 8 0 0 0 0 0 0 0 86 105 115 105 98 108 101 0 1 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 45 1 0 0 55 1 0 0 5 0 0 2 18 0 0 0 4 0 0 0 9 64 64 128 4 0 128 0 9 64 64 128 4 0 0 1 6 0 64 0 26 0 0 0 22 0 1 128 4 0 128 1 9 64 64 128 4 0 0 2 9 128 64 128 22 192 0 128 4 0 128 1 9 128 64 128 4 0 0 2 9 64 64 128 30 0 128 0 3 0 0 0 4 8 0 0 0 0 0 0 0 86 105 115 105 98 108 101 0 1 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 57 1 0 0 62 1 0 0 4 0 0 2 9 0 0 0 4 0 0 0 9 64 64 128 4 0 128 0 9 64 64 128 4 0 0 1 9 64 64 128 4 0 128 1 9 128 64 128 30 0 128 0 3 0 0 0 4 8 0 0 0 0 0 0 0 86 105 115 105 98 108 101 0 1 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 67 1 0 0 70 1 0 0 2 0 0 6 18 0 0 0 4 0 0 0 69 64 0 0 70 128 192 0 133 192 0 0 196 0 128 0 198 0 193 1 156 128 0 1 197 192 0 0 4 1 128 0 6 1 65 2 220 128 0 1 5 193 0 0 68 1 128 0 70 1 193 2 28 1 0 1 92 128 0 0 9 64 0 128 30 0 128 0 5 0 0 0 4 8 0 0 0 0 0 0 0 65 109 98 105 101 110 116 0 4 7 0 0 0 0 0 0 0 67 111 108 111 114 51 0 4 8 0 0 0 0 0 0 0 102 114 111 109 82 71 66 0 4 9 0 0 0 0 0 0 0 116 111 110 117 109 98 101 114 0 4 5 0 0 0 0 0 0 0 84 101 120 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 100 1 0 0 123 1 0 0 5 4 0 9 57 0 0 0 87 0 64 0 22 64 0 128 23 0 64 1 22 0 0 128 30 0 128 0 4 1 0 0 68 1 128 0 14 65 1 2 88 0 0 2 22 0 1 128 4 1 0 1 68 1 128 0 14 65 1 2 24 128 0 2 22 0 0 128 30 0 128 0 5 65 0 0 6 129 64 2 65 193 0 0 129 193 0 0 193 193 0 0 28 129 0 2 23 0 129 1 22 0 0 128 30 0 128 0 4 1 128 1 6 1 65 2 65 65 1 0 28 129 0 1 69 193 1 0 70 1 194 2 132 1 128 0 196 1 128 0 4 2 128 0 92 129 0 2 9 65 1 131 9 129 194 132 69 193 1 0 70 1 194 2 128 1 0 0 192 1 128 0 0 2 0 1 92 129 0 2 9 65 129 133 68 1 0 2 9 65 1 134 9 193 128 134 69 65 0 0 70 129 192 2 129 1 0 0 193 1 0 0 1 130 3 0 92 129 0 2 23 64 129 1 22 192 255 127 30 1 0 1 30 0 128 0 15 0 0 0 3 0 0 0 0 0 0 0 0 4 7 0 0 0 0 0 0 0 67 111 108 111 114 51 0 4 8 0 0 0 0 0 0 0 102 114 111 109 82 71 66 0 3 0 0 0 0 0 224 111 64 4 9 0 0 0 0 0 0 0 67 114 101 97 116 101 85 73 0 4 5 0 0 0 0 0 0 0 80 97 114 116 0 4 5 0 0 0 0 0 0 0 83 105 122 101 0 4 8 0 0 0 0 0 0 0 86 101 99 116 111 114 51 0 4 4 0 0 0 0 0 0 0 110 101 119 0 4 9 0 0 0 0 0 0 0 65 110 99 104 111 114 101 100 0 1 1 4 9 0 0 0 0 0 0 0 80 111 115 105 116 105 111 110 0 4 7 0 0 0 0 0 0 0 80 97 114 101 110 116 0 4 6 0 0 0 0 0 0 0 67 111 108 111 114 0 3 0 0 0 0 0 192 98 64 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 125 1 0 0 144 1 0 0 4 3 0 14 106 0 0 0 197 0 0 0 198 64 192 1 1 129 0 0 65 193 0 0 129 1 1 0 220 128 0 2 5 65 1 0 6 129 65 2 64 1 0 1 28 129 0 1 68 1 0 0 14 65 1 2 68 1 128 0 12 65 1 2 68 1 0 1 24 64 1 2 22 128 1 128 5 1 0 0 6 65 64 2 65 129 0 0 129 129 0 0 193 193 1 0 28 129 0 2 192 0 0 2 4 1 128 1 68 1 0 0 78 65 1 0 133 65 1 0 134 129 65 3 192 1 0 1 156 129 0 1 196 1 0 0 142 193 1 3 196 1 128 0 140 193 1 3 196 1 0 0 206 193 129 0 0 2 128 1 28 65 128 2 4 1 128 0 69 65 1 0 70 129 193 2 128 1 0 1 92 129 0 1 132 1 0 0 78 129 129 2 12 65 1 2 68 1 0 0 13 65 1 2 69 65 1 0 70 129 193 2 128 1 0 1 92 129 0 1 132 1 0 0 78 129 129 2 132 1 128 0 76 129 129 2 132 1 0 1 24 128 129 2 22 128 6 128 68 1 0 1 133 65 1 0 134 129 65 3 192 1 0 1 156 129 0 1 196 1 0 0 142 193 1 3 196 1 128 0 140 193 1 3 24 64 1 3 22 192 3 128 132 1 128 1 196 1 0 0 206 193 1 0 0 2 128 2 68 2 0 0 78 66 130 0 133 2 0 0 134 66 64 5 193 130 0 0 1 131 0 0 65 195 1 0 156 2 0 2 156 65 0 0 132 1 0 0 77 129 129 2 22 64 249 127 24 0 1 129 22 192 3 128 68 1 128 1 132 1 0 0 142 129 1 0 192 1 0 2 4 2 0 0 14 2 130 0 69 2 0 0 70 66 192 4 129 2 2 0 193 2 2 0 1 3 2 0 92 2 0 2 92 65 0 0 68 1 0 0 13 65 1 2 22 64 251 127 30 0 128 0 9 0 0 0 4 7 0 0 0 0 0 0 0 67 111 108 111 114 51 0 4 8 0 0 0 0 0 0 0 102 114 111 109 82 71 66 0 3 0 0 0 0 0 0 0 0 3 0 0 0 0 0 64 99 64 3 0 0 0 0 0 0 55 64 4 5 0 0 0 0 0 0 0 109 97 116 104 0 4 6 0 0 0 0 0 0 0 102 108 111 111 114 0 3 0 0 0 0 0 192 98 64 3 0 0 0 0 0 0 62 64 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 193 1 0 0 233 1 0 0 12 1 0 22 203 0 0 0 91 64 0 0 22 0 1 128 69 0 0 0 70 64 192 0 129 128 0 0 193 192 0 0 92 128 128 1 133 0 1 0 192 0 0 0 156 128 0 1 23 64 65 1 22 192 2 128 65 128 1 0 139 192 65 0 1 1 2 0 156 0 129 1 22 0 1 128 133 65 1 0 134 65 66 3 192 1 128 2 156 129 0 1 76 128 129 0 161 64 0 0 22 0 254 127 133 0 0 0 134 128 66 1 192 0 128 0 156 64 0 1 129 128 0 0 196 0 0 0 1 129 0 0 160 0 42 128 129 129 0 0 196 1 128 0 1 130 0 0 160 1 37 128 133 2 0 0 134 194 66 5 196 2 128 0 207 194 130 4 204 66 128 5 4 3 0 0 15 3 131 2 12 67 0 6 65 131 1 0 156 130 0 2 196 2 0 1 142 194 2 5 196 2 128 1 0 3 128 4 64 3 128 2 128 3 0 5 220 66 0 2 197 2 0 0 198 66 192 5 1 131 0 0 68 3 0 2 220 130 128 1 23 128 192 5 22 0 31 128 197 2 0 0 198 2 195 5 0 3 0 5 220 130 0 1 4 3 128 2 206 2 131 5 4 3 0 3 204 2 131 5 4 3 128 3 24 192 2 6 22 64 28 128 197 66 3 0 4 3 0 4 220 2 1 1 22 192 26 128 4 4 128 4 70 132 195 7 70 196 195 8 76 68 132 4 6 68 4 8 23 0 68 8 22 64 1 128 4 4 128 4 70 132 195 7 70 196 195 8 76 68 132 4 138 4 0 0 9 132 132 8 4 4 128 4 70 132 195 7 70 196 195 8 76 68 132 4 6 68 4 8 69 4 0 0 70 4 195 8 128 4 0 5 92 132 0 1 134 132 195 7 134 68 68 9 76 132 132 8 6 68 4 8 23 0 68 8 22 64 3 128 4 4 128 4 70 132 195 7 70 196 195 8 76 68 132 4 6 68 4 8 69 4 0 0 70 4 195 8 128 4 0 5 92 132 0 1 134 132 195 7 134 68 68 9 76 132 132 8 138 4 0 0 9 132 132 8 4 4 128 4 70 132 195 7 70 196 195 8 76 68 132 4 6 68 4 8 69 4 0 0 70 4 195 8 128 4 0 5 92 132 0 1 134 132 195 7 134 68 68 9 76 132 132 8 6 68 4 8 70 132 195 7 70 132 196 8 76 68 132 2 6 68 4 8 23 0 68 8 22 64 7 128 4 4 0 5 68 4 128 2 78 68 132 4 134 132 195 7 134 196 67 9 196 4 128 2 142 196 4 9 76 132 132 8 133 4 0 0 134 4 67 9 192 4 0 5 156 132 0 1 196 4 128 2 142 196 4 9 196 4 0 3 140 196 4 9 198 132 195 7 198 68 196 9 4 5 128 2 206 4 133 9 140 196 4 9 196 4 128 2 206 196 132 2 6 133 195 7 6 133 68 10 68 5 128 2 14 69 5 10 204 4 133 9 6 197 196 7 28 68 128 2 4 4 128 4 70 132 195 7 70 196 195 8 76 68 132 4 6 68 4 8 69 4 0 0 70 4 195 8 128 4 0 5 92 132 0 1 134 132 195 7 134 68 68 9 76 132 132 8 6 68 4 8 70 132 195 7 70 132 196 8 76 68 132 2 9 4 197 8 225 130 0 0 22 64 228 127 159 65 218 127 132 1 128 5 197 129 5 0 5 2 0 0 6 2 67 4 68 2 0 0 79 66 130 2 78 194 197 4 28 2 0 1 220 129 0 0 1 2 6 0 213 1 130 3 137 193 129 138 133 65 6 0 134 129 70 3 156 65 128 0 159 64 213 127 30 0 128 0 27 0 0 0 4 5 0 0 0 0 0 0 0 109 97 116 104 0 4 7 0 0 0 0 0 0 0 114 97 110 100 111 109 0 3 0 0 0 0 0 0 240 63 3 0 0 0 0 132 215 151 65 4 7 0 0 0 0 0 0 0 116 121 112 101 111 102 0 4 7 0 0 0 0 0 0 0 115 116 114 105 110 103 0 3 0 0 0 0 0 0 0 0 4 7 0 0 0 0 0 0 0 103 109 97 116 99 104 0 4 2 0 0 0 0 0 0 0 46 0 4 5 0 0 0 0 0 0 0 98 121 116 101 0 4 11 0 0 0 0 0 0 0 114 97 110 100 111 109 115 101 101 100 0 4 6 0 0 0 0 0 0 0 110 111 105 115 101 0 4 6 0 0 0 0 0 0 0 102 108 111 111 114 0 4 6 0 0 0 0 0 0 0 112 97 105 114 115 0 4 4 0 0 0 0 0 0 0 80 111 115 0 4 2 0 0 0 0 0 0 0 88 0 0 4 2 0 0 0 0 0 0 0 89 0 4 2 0 0 0 0 0 0 0 90 0 4 6 0 0 0 0 0 0 0 67 111 108 111 114 0 1 1 4 5 0 0 0 0 0 0 0 84 101 120 116 0 4 9 0 0 0 0 0 0 0 116 111 115 116 114 105 110 103 0 3 0 0 0 0 0 0 89 64 4 2 0 0 0 0 0 0 0 37 0 4 5 0 0 0 0 0 0 0 116 97 115 107 0 4 5 0 0 0 0 0 0 0 119 97 105 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 248 1 0 0 5 2 0 0 5 0 0 7 47 0 0 0 4 0 0 0 11 0 64 0 28 128 0 1 68 0 128 0 134 64 64 0 196 0 0 1 142 192 0 1 76 128 128 0 72 0 128 0 68 0 128 1 134 128 64 0 196 0 0 1 142 192 0 1 76 128 128 0 72 0 128 1 68 0 128 0 24 64 128 129 22 64 0 128 65 192 0 0 72 0 128 0 68 0 128 0 24 0 193 0 22 64 0 128 65 0 1 0 72 0 128 0 68 0 0 2 133 64 1 0 134 128 65 1 196 0 0 2 198 64 193 1 198 192 193 1 156 128 0 1 197 64 1 0 198 0 194 1 5 65 2 0 6 129 66 2 68 1 128 0 28 129 0 1 69 65 2 0 70 129 194 2 132 1 128 1 92 129 0 1 129 193 2 0 220 128 0 2 142 192 0 1 73 128 128 130 30 0 128 0 12 0 0 0 4 14 0 0 0 0 0 0 0 71 101 116 77 111 117 115 101 68 101 108 116 97 0 4 2 0 0 0 0 0 0 0 89 0 4 2 0 0 0 0 0 0 0 88 0 3 0 0 0 0 0 128 86 64 3 0 0 0 0 0 128 86 192 4 7 0 0 0 0 0 0 0 67 70 114 97 109 101 0 4 4 0 0 0 0 0 0 0 110 101 119 0 4 9 0 0 0 0 0 0 0 80 111 115 105 116 105 111 110 0 4 16 0 0 0 0 0 0 0 102 114 111 109 79 114 105 101 110 116 97 116 105 111 110 0 4 5 0 0 0 0 0 0 0 109 97 116 104 0 4 4 0 0 0 0 0 0 0 114 97 100 0 3 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 19 2 0 0 101 2 0 0 3 1 0 20 170 0 0 0 129 0 0 0 202 0 0 0 5 65 0 0 6 129 64 2 64 1 0 0 164 1 0 0 28 65 128 1 10 1 0 0 69 193 0 0 128 1 0 0 92 1 1 1 22 128 21 128 140 2 65 4 134 130 2 0 154 2 0 0 22 0 12 128 198 66 193 4 198 130 193 5 6 67 65 5 6 131 65 6 23 0 131 5 22 128 10 128 198 66 193 4 198 194 193 5 6 67 65 5 6 195 65 6 23 0 131 5 22 0 9 128 198 66 193 4 198 2 194 5 4 3 0 0 207 2 131 5 204 2 193 5 6 67 65 5 6 3 66 6 68 3 0 0 15 67 3 6 13 3 65 6 65 3 1 0 224 130 5 128 202 131 0 0 5 68 2 0 6 132 66 8 70 68 193 4 70 132 193 8 132 4 0 0 142 132 4 7 198 68 193 4 198 196 193 9 28 132 0 2 201 3 132 130 5 4 3 0 6 68 67 8 65 132 3 0 129 132 3 0 193 132 3 0 28 132 0 2 201 3 132 133 5 68 0 0 6 196 67 8 64 4 0 2 128 4 128 7 28 68 128 1 223 194 249 127 22 64 8 128 198 66 193 4 198 2 194 5 4 3 0 0 207 2 131 5 204 2 193 5 4 3 128 0 68 3 0 0 15 67 3 6 65 3 1 0 224 130 5 128 202 131 0 0 5 68 2 0 6 132 66 8 70 68 193 4 70 132 193 8 132 4 0 0 142 132 4 7 198 68 193 4 198 196 193 9 28 132 0 2 201 3 132 130 5 4 3 0 6 68 67 8 65 132 3 0 129 132 3 0 193 132 3 0 28 132 0 2 201 3 132 133 5 68 0 0 6 196 67 8 64 4 0 2 128 4 128 7 28 68 128 1 223 194 249 127 97 129 0 0 22 128 233 127 69 193 0 0 128 1 0 2 92 1 1 1 22 0 1 128 133 66 0 0 134 194 67 5 192 2 0 0 0 3 128 4 156 66 128 1 97 129 0 0 22 0 254 127 68 1 0 1 148 1 0 0 92 65 0 1 69 65 0 0 70 129 192 2 128 1 0 0 228 65 0 0 92 65 128 1 69 193 0 0 128 1 0 0 92 1 1 1 22 192 7 128 90 0 0 0 22 192 3 128 134 66 193 0 134 130 65 5 198 66 193 4 198 130 193 5 23 192 2 5 22 64 2 128 134 66 193 0 134 194 65 5 198 66 193 4 198 194 193 5 23 192 2 5 22 192 0 128 134 194 194 0 198 194 194 4 87 192 2 5 22 0 3 128 90 0 0 0 22 192 1 128 133 66 0 0 134 194 67 5 192 2 128 1 10 3 0 1 70 195 194 0 128 3 0 1 34 67 0 1 156 66 128 1 64 0 128 4 129 0 1 0 22 0 0 128 140 0 65 1 97 129 0 0 22 64 247 127 90 0 0 0 22 192 1 128 69 65 0 0 70 193 195 2 128 1 128 1 202 1 0 1 6 194 194 0 64 2 0 1 226 65 0 1 92 65 128 1 222 0 0 1 30 0 128 0 16 0 0 0 3 0 0 0 0 0 0 0 0 4 6 0 0 0 0 0 0 0 116 97 98 108 101 0 4 5 0 0 0 0 0 0 0 115 111 114 116 0 4 7 0 0 0 0 0 0 0 105 112 97 105 114 115 0 3 0 0 0 0 0 0 240 63 4 9 0 0 0 0 0 0 0 80 111 115 105 116 105 111 110 0 4 2 0 0 0 0 0 0 0 88 0 4 2 0 0 0 0 0 0 0 90 0 4 2 0 0 0 0 0 0 0 89 0 4 8 0 0 0 0 0 0 0 86 101 99 116 111 114 51 0 4 4 0 0 0 0 0 0 0 110 101 119 0 4 6 0 0 0 0 0 0 0 67 111 108 111 114 0 4 7 0 0 0 0 0 0 0 67 111 108 111 114 51 0 4 8 0 0 0 0 0 0 0 102 114 111 109 82 71 66 0 3 0 0 0 0 0 224 111 64 4 7 0 0 0 0 0 0 0 105 110 115 101 114 116 0 2 0 0 0 0 0 0 0 0 0 0 0 25 2 0 0 33 2 0 0 0 2 0 4 42 0 0 0 134 0 64 0 134 64 64 1 198 0 192 0 198 64 192 1 87 192 0 1 22 64 2 128 134 0 64 0 134 64 64 1 198 0 192 0 198 64 192 1 88 192 0 1 22 0 0 128 130 64 0 0 130 0 128 0 158 0 0 1 22 0 6 128 134 0 64 0 134 128 64 1 198 0 192 0 198 128 192 1 87 192 0 1 22 64 2 128 134 0 64 0 134 128 64 1 198 0 192 0 198 128 192 1 88 192 0 1 22 0 0 128 130 64 0 0 130 0 128 0 158 0 0 1 22 0 2 128 134 0 64 0 134 192 64 1 198 0 192 0 198 192 192 1 88 192 0 1 22 0 0 128 130 64 0 0 130 0 128 0 158 0 0 1 30 0 128 0 4 0 0 0 4 9 0 0 0 0 0 0 0 80 111 115 105 116 105 111 110 0 4 2 0 0 0 0 0 0 0 88 0 4 2 0 0 0 0 0 0 0 90 0 4 2 0 0 0 0 0 0 0 89 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 70 2 0 0 78 2 0 0 0 2 0 4 42 0 0 0 134 0 64 0 134 64 64 1 198 0 192 0 198 64 192 1 87 192 0 1 22 64 2 128 134 0 64 0 134 64 64 1 198 0 192 0 198 64 192 1 88 192 0 1 22 0 0 128 130 64 0 0 130 0 128 0 158 0 0 1 22 0 6 128 134 0 64 0 134 128 64 1 198 0 192 0 198 128 192 1 87 192 0 1 22 64 2 128 134 0 64 0 134 128 64 1 198 0 192 0 198 128 192 1 88 192 0 1 22 0 0 128 130 64 0 0 130 0 128 0 158 0 0 1 22 0 2 128 134 0 64 0 134 192 64 1 198 0 192 0 198 192 192 1 88 192 0 1 22 0 0 128 130 64 0 0 130 0 128 0 158 0 0 1 30 0 128 0 4 0 0 0 4 9 0 0 0 0 0 0 0 80 111 115 105 116 105 111 110 0 4 2 0 0 0 0 0 0 0 88 0 4 2 0 0 0 0 0 0 0 90 0 4 2 0 0 0 0 0 0 0 89 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 103 2 0 0 128 2 0 0 5 1 0 20 47 0 0 0 65 0 0 0 129 0 0 0 193 0 0 0 4 1 0 0 84 1 0 0 28 65 0 1 5 65 0 0 64 1 0 0 28 1 1 1 22 64 8 128 70 2 64 4 133 130 0 0 198 194 64 4 156 130 0 1 193 2 0 0 0 3 0 5 65 3 0 0 224 2 6 128 196 3 128 0 4 4 0 1 14 4 132 0 68 4 0 1 78 68 4 1 132 4 0 1 142 132 132 1 192 4 128 4 220 67 128 2 140 0 64 1 196 3 128 1 4 4 0 1 207 3 132 7 204 3 192 7 23 192 3 1 22 64 0 128 129 0 0 0 76 0 192 0 196 3 0 2 204 3 192 7 23 192 131 0 22 128 0 128 129 0 0 0 65 0 0 0 204 0 192 1 223 66 249 127 33 129 0 0 22 192 246 127 30 0 128 0 4 0 0 0 3 0 0 0 0 0 0 240 63 4 7 0 0 0 0 0 0 0 105 112 97 105 114 115 0 4 9 0 0 0 0 0 0 0 116 111 110 117 109 98 101 114 0 3 0 0 0 0 0 0 0 64 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 130 2 0 0 141 2 0 0 4 1 0 14 44 0 0 0 74 0 0 0 133 0 0 0 192 0 0 0 156 0 1 1 22 0 4 128 197 65 0 0 198 129 192 3 4 2 0 0 70 194 64 3 220 129 128 1 87 0 193 3 22 64 2 128 5 66 0 0 6 66 65 4 64 2 128 0 133 130 1 0 134 194 65 5 193 2 2 0 0 3 128 3 70 67 66 3 156 2 0 2 28 66 0 0 161 128 0 0 22 0 251 127 133 64 0 0 134 128 66 1 202 0 128 1 4 1 128 0 68 1 0 1 132 1 128 1 226 64 128 1 1 193 2 0 156 128 128 1 193 0 3 0 149 192 0 1 192 0 0 1 5 65 0 0 6 129 66 2 64 1 128 0 129 65 3 0 28 129 128 1 149 0 129 1 158 0 0 1 30 0 128 0 14 0 0 0 4 7 0 0 0 0 0 0 0 105 112 97 105 114 115 0 4 6 0 0 0 0 0 0 0 116 97 98 108 101 0 4 5 0 0 0 0 0 0 0 102 105 110 100 0 3 0 0 0 0 0 0 240 63 0 4 7 0 0 0 0 0 0 0 105 110 115 101 114 116 0 4 7 0 0 0 0 0 0 0 115 116 114 105 110 103 0 4 7 0 0 0 0 0 0 0 102 111 114 109 97 116 0 4 6 0 0 0 0 0 0 0 37 100 124 37 100 0 3 0 0 0 0 0 0 0 64 4 7 0 0 0 0 0 0 0 99 111 110 99 97 116 0 4 2 0 0 0 0 0 0 0 46 0 4 2 0 0 0 0 0 0 0 44 0 4 2 0 0 0 0 0 0 0 126 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 143 2 0 0 159 2 0 0 4 1 0 16 50 0 0 0 74 0 0 0 139 0 64 0 1 65 0 0 156 128 128 1 134 128 64 1 139 0 64 1 1 193 0 0 156 128 128 1 197 0 1 0 6 129 64 1 220 128 0 1 200 0 0 0 197 0 1 0 6 65 65 1 220 128 0 1 200 0 128 0 197 0 1 0 6 129 65 1 220 128 0 1 200 0 0 1 203 0 64 0 65 65 0 0 220 128 128 1 198 64 193 1 203 0 192 1 65 193 1 0 220 128 128 1 5 1 2 0 64 1 128 1 28 1 1 1 22 128 3 128 75 2 64 4 193 66 2 0 92 130 128 1 133 2 1 0 198 130 192 4 156 130 0 1 197 130 2 0 198 194 194 5 0 3 128 0 74 3 0 1 132 3 128 1 134 131 2 7 198 67 193 4 98 67 0 1 220 66 128 1 33 129 0 0 22 128 251 127 94 0 0 1 30 0 128 0 12 0 0 0 4 6 0 0 0 0 0 0 0 115 112 108 105 116 0 4 2 0 0 0 0 0 0 0 44 0 3 0 0 0 0 0 0 240 63 4 2 0 0 0 0 0 0 0 46 0 4 9 0 0 0 0 0 0 0 116 111 110 117 109 98 101 114 0 3 0 0 0 0 0 0 0 64 3 0 0 0 0 0 0 8 64 4 2 0 0 0 0 0 0 0 126 0 4 7 0 0 0 0 0 0 0 105 112 97 105 114 115 0 4 2 0 0 0 0 0 0 0 124 0 4 6 0 0 0 0 0 0 0 116 97 98 108 101 0 4 7 0 0 0 0 0 0 0 105 110 115 101 114 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 161 2 0 0 171 2 0 0 4 1 0 8 67 0 0 0 68 0 0 0 70 0 192 0 132 0 0 0 134 64 64 1 156 128 128 0 193 128 0 0 0 1 0 0 65 193 0 0 149 64 1 1 92 128 0 1 90 0 0 0 22 64 2 128 68 0 0 0 70 0 193 0 132 0 0 0 134 64 64 1 156 128 128 0 193 128 0 0 0 1 0 0 65 193 0 0 149 64 1 1 92 64 0 1 68 0 0 0 70 64 193 0 132 0 0 0 134 64 64 1 156 128 128 0 193 128 0 0 0 1 0 0 65 193 0 0 149 64 1 1 195 0 128 1 1 129 1 0 92 64 0 2 68 0 128 0 75 192 193 0 92 128 0 1 133 0 2 0 193 64 2 0 5 129 2 0 84 1 128 0 28 129 0 1 65 193 2 0 213 64 129 1 156 64 0 1 133 0 3 0 134 64 67 1 156 64 128 0 132 0 0 1 196 0 128 1 0 1 128 0 220 0 0 1 156 128 0 0 196 0 0 0 198 128 195 1 4 1 0 0 6 65 64 2 28 129 128 0 65 129 0 0 128 1 0 0 193 193 0 0 21 193 1 2 64 1 0 1 131 1 0 3 194 1 128 0 220 64 128 2 30 0 128 0 15 0 0 0 4 11 0 0 0 0 0 0 0 70 105 108 101 69 120 105 115 116 115 0 4 17 0 0 0 0 0 0 0 71 101 116 79 83 68 114 105 118 101 76 101 116 116 101 114 0 4 35 0 0 0 0 0 0 0 58 47 83 121 115 116 101 109 47 65 112 112 68 97 116 97 47 66 117 105 108 100 66 114 101 97 107 47 115 97 118 101 115 47 0 4 5 0 0 0 0 0 0 0 46 100 97 116 0 4 13 0 0 0 0 0 0 0 68 101 108 101 116 101 79 98 106 101 99 116 0 4 11 0 0 0 0 0 0 0 67 114 101 97 116 101 70 105 108 101 0 4 8 0 0 0 0 0 0 0 82 45 87 45 68 45 65 0 4 12 0 0 0 0 0 0 0 71 101 116 67 104 105 108 100 114 101 110 0 4 6 0 0 0 0 0 0 0 112 114 105 110 116 0 4 8 0 0 0 0 0 0 0 115 97 118 105 110 103 32 0 4 9 0 0 0 0 0 0 0 116 111 115 116 114 105 110 103 0 4 7 0 0 0 0 0 0 0 32 112 97 114 116 115 0 4 5 0 0 0 0 0 0 0 116 97 115 107 0 4 5 0 0 0 0 0 0 0 119 97 105 116 0 4 10 0 0 0 0 0 0 0 87 114 105 116 101 70 105 108 101 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 172 2 0 0 175 2 0 0 2 1 0 5 16 0 0 0 68 0 0 0 70 0 192 0 132 0 0 0 134 64 64 1 156 128 128 0 193 128 0 0 0 1 0 0 149 0 1 1 92 128 0 1 70 192 192 0 133 0 1 0 196 0 128 0 0 1 128 0 220 0 0 1 156 64 0 0 30 0 128 0 5 0 0 0 4 8 0 0 0 0 0 0 0 71 101 116 70 105 108 101 0 4 17 0 0 0 0 0 0 0 71 101 116 79 83 68 114 105 118 101 76 101 116 116 101 114 0 4 35 0 0 0 0 0 0 0 58 47 83 121 115 116 101 109 47 65 112 112 68 97 116 97 47 66 117 105 108 100 66 114 101 97 107 47 115 97 118 101 115 47 0 4 5 0 0 0 0 0 0 0 68 97 116 97 0 4 11 0 0 0 0 0 0 0 86 82 76 69 100 101 99 111 100 101 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 191 2 0 0 196 2 0 0 3 0 0 5 17 0 0 0 4 0 0 0 11 0 64 0 132 0 128 0 134 64 64 1 134 128 64 1 196 0 128 0 198 64 192 1 198 192 192 1 4 1 0 1 206 0 129 1 28 128 0 2 26 0 0 0 22 128 0 128 70 0 65 0 75 64 193 0 92 64 0 1 30 0 128 0 6 0 0 0 4 8 0 0 0 0 0 0 0 82 97 121 99 97 115 116 0 4 7 0 0 0 0 0 0 0 67 70 114 97 109 101 0 4 9 0 0 0 0 0 0 0 80 111 115 105 116 105 111 110 0 4 11 0 0 0 0 0 0 0 76 111 111 107 86 101 99 116 111 114 0 4 9 0 0 0 0 0 0 0 73 110 115 116 97 110 99 101 0 4 8 0 0 0 0 0 0 0 68 101 115 116 114 111 121 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 198 2 0 0 205 2 0 0 5 0 0 11 43 0 0 0 4 0 0 0 11 0 64 0 132 0 128 0 134 64 64 1 134 128 64 1 196 0 128 0 198 64 192 1 198 192 192 1 4 1 0 1 206 0 129 1 28 128 0 2 26 0 0 0 22 0 7 128 69 0 1 0 70 64 193 0 134 128 65 0 134 192 65 1 196 0 128 1 142 192 0 1 198 128 65 0 198 0 194 1 4 1 128 1 206 0 129 1 6 129 65 0 6 65 66 2 68 1 128 1 14 65 1 2 92 128 0 2 134 128 66 0 134 128 64 1 140 64 0 1 196 0 0 2 6 193 65 1 70 1 66 1 134 65 66 1 197 193 2 0 198 1 195 3 1 66 3 0 65 130 3 0 129 194 3 0 220 1 0 2 220 64 0 0 30 0 128 0 16 0 0 0 4 8 0 0 0 0 0 0 0 82 97 121 99 97 115 116 0 4 7 0 0 0 0 0 0 0 67 70 114 97 109 101 0 4 9 0 0 0 0 0 0 0 80 111 115 105 116 105 111 110 0 4 11 0 0 0 0 0 0 0 76 111 111 107 86 101 99 116 111 114 0 4 8 0 0 0 0 0 0 0 86 101 99 116 111 114 51 0 4 4 0 0 0 0 0 0 0 110 101 119 0 4 7 0 0 0 0 0 0 0 78 111 114 109 97 108 0 4 2 0 0 0 0 0 0 0 88 0 4 2 0 0 0 0 0 0 0 89 0 4 2 0 0 0 0 0 0 0 90 0 4 9 0 0 0 0 0 0 0 73 110 115 116 97 110 99 101 0 4 7 0 0 0 0 0 0 0 67 111 108 111 114 51 0 4 8 0 0 0 0 0 0 0 102 114 111 109 82 71 66 0 3 0 0 0 0 0 128 100 64 3 0 0 0 0 0 0 93 64 3 0 0 0 0 0 64 82 64 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 207 2 0 0 214 2 0 0 2 0 0 2 18 0 0 0 4 0 0 0 6 0 64 0 69 64 0 0 70 0 192 0 70 128 192 0 23 64 0 0 22 192 1 128 4 0 0 0 69 64 0 0 70 0 192 0 70 192 192 0 9 64 0 128 4 0 0 0 9 64 65 130 22 64 0 128 4 0 128 0 28 64 128 0 30 0 128 0 6 0 0 0 4 14 0 0 0 0 0 0 0 77 111 117 115 101 66 101 104 97 118 105 111 114 0 4 5 0 0 0 0 0 0 0 69 110 117 109 0 4 8 0 0 0 0 0 0 0 68 101 102 97 117 108 116 0 4 20 0 0 0 0 0 0 0 76 111 99 107 67 117 114 114 101 110 116 80 111 115 105 116 105 111 110 0 4 17 0 0 0 0 0 0 0 77 111 117 115 101 73 99 111 110 69 110 97 98 108 101 100 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 216 2 0 0 221 2 0 0 2 0 0 2 11 0 0 0 4 0 0 0 6 0 64 0 69 64 0 0 70 0 192 0 70 128 192 0 23 64 0 0 22 0 0 128 30 0 128 0 4 0 128 0 28 64 128 0 30 0 128 0 3 0 0 0 4 14 0 0 0 0 0 0 0 77 111 117 115 101 66 101 104 97 118 105 111 114 0 4 5 0 0 0 0 0 0 0 69 110 117 109 0 4 8 0 0 0 0 0 0 0 68 101 102 97 117 108 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 223 2 0 0 228 2 0 0 2 0 0 2 11 0 0 0 4 0 0 0 6 0 64 0 69 64 0 0 70 0 192 0 70 128 192 0 23 64 0 0 22 0 0 128 30 0 128 0 4 0 128 0 28 64 128 0 30 0 128 0 3 0 0 0 4 14 0 0 0 0 0 0 0 77 111 117 115 101 66 101 104 97 118 105 111 114 0 4 5 0 0 0 0 0 0 0 69 110 117 109 0 4 8 0 0 0 0 0 0 0 68 101 102 97 117 108 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 230 2 0 0 235 2 0 0 2 0 0 2 11 0 0 0 4 0 0 0 6 0 64 0 69 64 0 0 70 0 192 0 70 128 192 0 23 64 0 0 22 0 0 128 30 0 128 0 4 0 128 0 28 64 128 0 30 0 128 0 3 0 0 0 4 14 0 0 0 0 0 0 0 77 111 117 115 101 66 101 104 97 118 105 111 114 0 4 5 0 0 0 0 0 0 0 69 110 117 109 0 4 8 0 0 0 0 0 0 0 68 101 102 97 117 108 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 237 2 0 0 245 2 0 0 2 1 0 5 17 0 0 0 68 0 0 0 70 0 192 0 129 64 0 0 92 128 0 1 129 192 0 0 192 0 0 0 149 192 0 1 73 128 0 129 132 0 128 0 139 0 65 1 0 1 128 0 156 64 128 1 133 64 1 0 228 0 0 0 0 0 128 0 156 64 0 1 30 0 128 0 6 0 0 0 4 9 0 0 0 0 0 0 0 67 114 101 97 116 101 85 73 0 4 6 0 0 0 0 0 0 0 83 111 117 110 100 0 4 8 0 0 0 0 0 0 0 83 111 117 110 100 73 100 0 4 14 0 0 0 0 0 0 0 114 98 120 97 115 115 101 116 105 100 58 47 47 0 4 15 0 0 0 0 0 0 0 80 108 97 121 76 111 99 97 108 83 111 117 110 100 0 4 6 0 0 0 0 0 0 0 115 112 97 119 110 0 1 0 0 0 0 0 0 0 0 0 0 0 241 2 0 0 244 2 0 0 1 0 0 2 8 0 0 0 4 0 0 0 6 0 64 0 11 64 64 0 28 64 0 1 4 0 0 0 11 128 64 0 28 64 0 1 30 0 128 0 3 0 0 0 4 6 0 0 0 0 0 0 0 69 110 100 101 100 0 4 5 0 0 0 0 0 0 0 87 97 105 116 0 4 8 0 0 0 0 0 0 0 68 101 115 116 114 111 121 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 247 2 0 0 11 3 0 0 6 2 0 8 77 0 0 0 134 0 64 0 197 64 0 0 198 0 192 1 198 128 192 1 23 192 0 1 22 64 8 128 132 0 0 0 134 192 64 1 23 0 65 1 22 64 7 128 132 0 128 0 134 64 65 1 197 64 0 0 198 64 193 1 198 128 193 1 23 192 0 1 22 192 2 128 132 0 128 0 197 64 0 0 198 64 193 1 198 192 193 1 137 192 128 130 132 0 128 0 137 64 66 132 132 0 0 1 137 64 194 129 132 0 128 1 137 0 193 129 22 128 2 128 132 0 128 0 197 64 0 0 198 64 193 1 198 128 193 1 137 192 128 130 132 0 128 0 137 0 65 132 132 0 128 1 137 64 194 129 132 0 0 1 137 0 193 129 134 0 64 0 197 64 0 0 198 0 192 1 198 128 194 1 23 192 0 1 22 128 4 128 90 64 0 0 22 0 4 128 132 0 0 2 197 192 2 0 198 0 195 1 5 65 3 0 6 1 67 2 68 1 0 2 70 193 194 2 70 129 195 2 70 193 195 2 129 1 4 0 196 1 0 2 198 193 194 3 198 129 195 3 198 65 196 3 28 1 0 2 220 128 0 0 137 192 128 133 134 0 64 0 197 64 0 0 198 0 192 1 198 128 196 1 23 192 0 1 22 0 1 128 90 64 0 0 22 128 0 128 132 0 128 2 193 192 4 0 156 64 0 1 30 0 128 0 20 0 0 0 4 8 0 0 0 0 0 0 0 75 101 121 67 111 100 101 0 4 5 0 0 0 0 0 0 0 69 110 117 109 0 4 4 0 0 0 0 0 0 0 84 97 98 0 4 8 0 0 0 0 0 0 0 86 105 115 105 98 108 101 0 1 1 4 14 0 0 0 0 0 0 0 77 111 117 115 101 66 101 104 97 118 105 111 114 0 4 8 0 0 0 0 0 0 0 68 101 102 97 117 108 116 0 4 20 0 0 0 0 0 0 0 76 111 99 107 67 117 114 114 101 110 116 80 111 115 105 116 105 111 110 0 4 17 0 0 0 0 0 0 0 77 111 117 115 101 73 99 111 110 69 110 97 98 108 101 100 0 1 0 4 2 0 0 0 0 0 0 0 82 0 4 7 0 0 0 0 0 0 0 67 70 114 97 109 101 0 4 4 0 0 0 0 0 0 0 110 101 119 0 4 8 0 0 0 0 0 0 0 86 101 99 116 111 114 51 0 4 9 0 0 0 0 0 0 0 80 111 115 105 116 105 111 110 0 4 2 0 0 0 0 0 0 0 88 0 3 0 0 0 0 0 0 94 64 4 2 0 0 0 0 0 0 0 90 0 4 2 0 0 0 0 0 0 0 69 0 3 64 250 4 28 230 60 219 66 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 13 3 0 0 18 3 0 0 3 0 0 2 12 0 0 0 4 0 0 0 69 64 0 0 70 0 192 0 70 128 192 0 9 64 0 128 4 0 0 0 9 0 193 129 4 0 128 0 9 128 193 130 4 0 0 1 9 0 193 130 30 0 128 0 7 0 0 0 4 14 0 0 0 0 0 0 0 77 111 117 115 101 66 101 104 97 118 105 111 114 0 4 5 0 0 0 0 0 0 0 69 110 117 109 0 4 20 0 0 0 0 0 0 0 76 111 99 107 67 117 114 114 101 110 116 80 111 115 105 116 105 111 110 0 4 17 0 0 0 0 0 0 0 77 111 117 115 101 73 99 111 110 69 110 97 98 108 101 100 0 1 0 4 8 0 0 0 0 0 0 0 86 105 115 105 98 108 101 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 20 3 0 0 27 3 0 0 7 0 0 3 19 0 0 0 4 0 0 0 11 0 64 0 28 64 0 1 4 0 128 0 6 64 64 0 65 128 0 0 132 0 0 1 28 128 128 1 8 0 0 0 4 0 128 1 11 192 64 0 28 64 0 1 4 0 0 2 9 64 65 130 4 0 128 2 9 64 65 130 4 0 0 3 9 128 65 130 30 0 128 0 7 0 0 0 4 8 0 0 0 0 0 0 0 68 101 115 116 114 111 121 0 4 9 0 0 0 0 0 0 0 67 114 101 97 116 101 85 73 0 4 7 0 0 0 0 0 0 0 70 111 108 100 101 114 0 4 11 0 0 0 0 0 0 0 68 105 115 99 111 110 110 101 99 116 0 4 8 0 0 0 0 0 0 0 86 105 115 105 98 108 101 0 1 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 42 3 0 0 53 3 0 0 1 1 0 8 24 0 0 0 74 0 0 0 133 0 0 0 134 64 64 1 156 128 128 0 196 0 0 0 203 128 192 1 70 193 64 0 134 1 65 0 192 1 0 1 220 128 128 2 218 0 0 0 22 192 1 128 11 65 65 1 134 129 193 1 28 65 128 1 5 193 1 0 6 1 66 2 64 1 128 0 128 1 128 1 28 65 128 1 218 64 0 0 22 64 251 127 94 0 0 1 30 0 128 0 9 0 0 0 4 14 0 0 0 0 0 0 0 82 97 121 99 97 115 116 80 97 114 97 109 115 0 4 4 0 0 0 0 0 0 0 110 101 119 0 4 8 0 0 0 0 0 0 0 82 97 121 99 97 115 116 0 4 7 0 0 0 0 0 0 0 79 114 105 103 105 110 0 4 10 0 0 0 0 0 0 0 68 105 114 101 99 116 105 111 110 0 4 12 0 0 0 0 0 0 0 65 100 100 84 111 70 105 108 116 101 114 0 4 9 0 0 0 0 0 0 0 73 110 115 116 97 110 99 101 0 4 6 0 0 0 0 0 0 0 116 97 98 108 101 0 4 7 0 0 0 0 0 0 0 105 110 115 101 114 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 55 3 0 0 83 3 0 0 3 1 0 12 92 0 0 0 68 0 0 0 133 0 0 0 134 64 64 1 197 128 0 0 198 64 192 1 4 1 128 0 6 193 64 2 6 1 65 2 6 65 65 2 68 1 128 0 70 193 192 2 70 1 193 2 70 129 193 2 77 193 193 2 132 1 128 0 134 193 64 3 134 1 65 3 134 1 66 3 220 128 0 2 5 129 0 0 6 65 64 2 70 65 65 0 134 65 65 0 24 128 129 132 22 128 0 128 132 1 0 1 154 65 0 0 22 192 1 128 134 65 65 0 24 64 66 3 22 192 0 128 132 1 0 1 146 1 0 3 154 65 0 0 22 0 0 128 129 65 2 0 76 129 129 2 134 129 65 0 198 1 66 0 6 2 66 0 24 0 130 132 22 128 0 128 4 2 0 1 26 66 0 0 22 192 1 128 6 2 66 0 24 64 66 4 22 192 0 128 4 2 0 1 18 2 0 4 26 66 0 0 22 0 0 128 1 66 2 0 204 1 130 3 28 1 0 2 156 0 0 0 92 128 0 0 148 0 128 0 24 128 128 132 22 64 7 128 133 128 0 0 134 64 64 1 193 64 2 0 1 65 2 0 65 65 2 0 156 128 0 2 197 128 2 0 0 1 128 0 220 0 1 1 22 0 4 128 6 194 194 3 18 2 0 4 70 194 194 3 78 66 2 0 70 2 195 4 14 66 2 4 77 2 2 0 132 2 128 0 134 194 64 5 134 2 65 5 140 66 2 5 196 2 128 0 198 194 192 5 198 2 193 5 205 194 2 5 140 192 2 1 22 64 0 128 225 128 0 0 22 0 251 127 158 0 0 1 30 0 0 1 30 0 128 0 13 0 0 0 4 4 0 0 0 0 0 0 0 82 97 121 0 4 4 0 0 0 0 0 0 0 110 101 119 0 4 8 0 0 0 0 0 0 0 86 101 99 116 111 114 51 0 4 7 0 0 0 0 0 0 0 67 70 114 97 109 101 0 4 9 0 0 0 0 0 0 0 80 111 115 105 116 105 111 110 0 4 2 0 0 0 0 0 0 0 88 0 4 2 0 0 0 0 0 0 0 89 0 3 0 0 0 0 0 0 240 63 4 2 0 0 0 0 0 0 0 90 0 3 0 0 0 0 0 0 0 0 4 6 0 0 0 0 0 0 0 112 97 105 114 115 0 4 7 0 0 0 0 0 0 0 78 111 114 109 97 108 0 4 10 0 0 0 0 0 0 0 77 97 103 110 105 116 117 100 101 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 85 3 0 0 131 3 0 0 15 0 0 4 23 0 0 0 4 0 0 0 6 0 64 0 65 64 0 0 28 128 0 1 70 128 64 0 75 192 192 0 228 0 0 0 4 0 0 1 4 0 128 1 4 0 0 2 4 0 128 2 4 0 0 3 4 0 128 3 4 0 0 4 4 0 128 4 4 0 0 5 4 0 128 5 4 0 0 6 4 0 128 6 4 0 0 7 92 128 128 1 72 0 128 0 30 0 128 0 4 0 0 0 4 11 0 0 0 0 0 0 0 71 101 116 83 101 114 118 105 99 101 0 4 11 0 0 0 0 0 0 0 82 117 110 83 101 114 118 105 99 101 0 4 14 0 0 0 0 0 0 0 82 101 110 100 101 114 83 116 101 112 112 101 100 0 4 8 0 0 0 0 0 0 0 67 111 110 110 101 99 116 0 1 0 0 0 0 0 0 0 0 0 0 0 87 3 0 0 130 3 0 0 13 1 0 10 13 1 0 0 68 0 0 0 70 0 192 0 133 64 0 0 134 0 64 1 134 128 64 1 23 128 128 0 22 0 0 128 30 0 128 0 68 0 0 0 75 192 192 0 197 64 0 0 198 0 193 1 198 64 193 1 92 128 128 1 90 0 0 0 22 192 6 128 68 0 128 0 70 128 193 0 70 192 193 0 75 0 194 0 197 64 2 0 198 128 194 1 1 193 2 0 65 1 3 0 129 193 2 0 220 0 0 2 92 128 0 0 82 0 128 0 132 0 128 0 196 0 128 0 198 128 193 1 4 1 0 1 69 65 2 0 70 129 194 2 134 65 195 0 193 193 2 0 6 130 195 0 92 129 0 2 132 1 128 1 142 1 0 3 78 129 129 2 28 129 0 1 204 0 129 1 137 192 0 131 68 0 0 0 75 192 192 0 197 64 0 0 198 0 193 1 198 192 195 1 92 128 128 1 90 0 0 0 22 0 7 128 68 0 128 0 70 128 193 0 70 192 193 0 75 0 194 0 197 64 2 0 198 128 194 1 1 193 2 0 65 1 3 0 129 193 2 0 220 0 0 2 92 128 0 0 82 0 128 0 132 0 128 0 196 0 128 0 198 128 193 1 4 1 0 1 69 65 2 0 70 129 194 2 134 65 195 0 193 193 2 0 6 130 195 0 92 129 0 2 132 1 128 1 142 1 0 3 146 1 0 3 78 129 129 2 28 129 0 1 204 0 129 1 137 192 0 131 68 0 0 0 75 192 192 0 197 64 0 0 198 0 193 1 198 0 196 1 92 128 128 1 90 0 0 0 22 0 7 128 68 0 128 0 70 128 193 0 133 128 1 0 134 64 68 1 193 192 2 0 5 129 4 0 6 193 68 2 65 1 5 0 28 129 0 1 65 193 2 0 156 128 0 2 78 128 128 0 70 64 197 0 132 0 128 0 196 0 128 0 198 128 193 1 4 1 0 1 69 65 2 0 70 129 194 2 134 65 195 0 193 193 2 0 6 130 195 0 92 129 0 2 132 1 128 1 142 1 0 3 78 129 129 2 28 129 0 1 204 0 129 1 137 192 0 131 68 0 0 0 75 192 192 0 197 64 0 0 198 0 193 1 198 128 197 1 92 128 128 1 90 0 0 0 22 0 7 128 68 0 128 0 70 128 193 0 133 128 1 0 134 64 68 1 193 192 2 0 5 129 4 0 6 193 68 2 65 193 5 0 28 129 0 1 65 193 2 0 156 128 0 2 78 128 128 0 70 64 197 0 132 0 128 0 196 0 128 0 198 128 193 1 4 1 0 1 69 65 2 0 70 129 194 2 134 65 195 0 193 193 2 0 6 130 195 0 92 129 0 2 132 1 128 1 142 1 0 3 78 129 129 2 28 129 0 1 204 0 129 1 137 192 0 131 68 0 0 2 75 0 198 0 196 0 128 0 198 128 193 1 198 64 198 1 5 65 2 0 6 129 66 2 65 193 2 0 132 1 128 2 196 1 0 3 140 193 1 3 146 1 0 3 193 193 2 0 28 1 0 2 92 128 0 0 132 0 0 0 139 192 64 1 5 65 0 0 6 1 65 2 6 129 70 2 156 128 128 1 154 0 0 0 22 64 1 128 90 0 0 0 22 192 0 128 132 0 0 4 142 128 128 141 136 0 128 3 66 0 0 0 132 0 128 3 196 0 128 4 206 0 128 1 140 192 0 1 136 0 128 3 132 0 128 3 196 0 0 5 209 0 128 1 142 192 0 1 136 0 128 3 90 64 0 0 22 0 3 128 132 0 128 0 196 0 128 0 198 128 193 1 5 65 2 0 6 129 66 2 65 193 2 0 132 1 128 3 142 1 0 3 193 193 2 0 28 129 0 2 204 0 129 1 137 192 0 131 22 128 4 128 129 192 2 0 136 0 128 3 132 0 128 0 196 0 128 0 198 128 193 1 6 65 198 0 69 65 2 0 70 129 194 2 129 193 2 0 196 1 0 3 1 194 2 0 92 129 0 2 12 65 1 2 68 1 128 0 70 129 193 2 70 65 198 2 13 65 1 2 204 0 129 1 137 192 0 131 132 0 128 5 197 128 4 0 198 64 199 1 15 1 0 134 220 128 0 1 1 129 7 0 213 0 129 1 137 192 0 142 132 0 0 6 197 128 4 0 198 64 199 1 4 1 128 0 6 129 65 2 6 65 70 2 6 65 67 2 68 1 0 4 15 65 1 2 220 128 0 1 1 193 7 0 69 129 4 0 70 65 199 2 132 1 128 0 134 129 65 3 134 65 70 3 134 1 72 3 196 1 0 4 143 193 1 3 92 129 0 1 129 193 7 0 197 129 4 0 198 65 199 3 4 2 128 0 6 130 65 4 6 66 70 4 6 130 67 4 68 2 0 4 15 66 2 4 220 129 0 1 213 192 129 1 137 192 0 142 30 0 128 0 33 0 0 0 4 14 0 0 0 0 0 0 0 77 111 117 115 101 66 101 104 97 118 105 111 114 0 4 5 0 0 0 0 0 0 0 69 110 117 109 0 4 8 0 0 0 0 0 0 0 68 101 102 97 117 108 116 0 4 10 0 0 0 0 0 0 0 73 115 75 101 121 68 111 119 110 0 4 8 0 0 0 0 0 0 0 75 101 121 67 111 100 101 0 4 2 0 0 0 0 0 0 0 87 0 4 7 0 0 0 0 0 0 0 67 70 114 97 109 101 0 4 12 0 0 0 0 0 0 0 82 105 103 104 116 86 101 99 116 111 114 0 4 6 0 0 0 0 0 0 0 67 114 111 115 115 0 4 8 0 0 0 0 0 0 0 86 101 99 116 111 114 51 0 4 4 0 0 0 0 0 0 0 110 101 119 0 3 0 0 0 0 0 0 0 0 3 0 0 0 0 0 0 240 63 4 2 0 0 0 0 0 0 0 88 0 4 2 0 0 0 0 0 0 0 90 0 4 2 0 0 0 0 0 0 0 83 0 4 2 0 0 0 0 0 0 0 65 0 4 7 0 0 0 0 0 0 0 65 110 103 108 101 115 0 4 5 0 0 0 0 0 0 0 109 97 116 104 0 4 4 0 0 0 0 0 0 0 114 97 100 0 3 0 0 0 0 0 128 86 64 4 11 0 0 0 0 0 0 0 76 111 111 107 86 101 99 116 111 114 0 4 2 0 0 0 0 0 0 0 68 0 3 0 0 0 0 0 128 86 192 4 8 0 0 0 0 0 0 0 82 97 121 99 97 115 116 0 4 9 0 0 0 0 0 0 0 80 111 115 105 116 105 111 110 0 4 6 0 0 0 0 0 0 0 83 112 97 99 101 0 3 0 0 0 0 0 0 16 64 4 5 0 0 0 0 0 0 0 84 101 120 116 0 4 6 0 0 0 0 0 0 0 102 108 111 111 114 0 4 5 0 0 0 0 0 0 0 32 70 80 83 0 4 2 0 0 0 0 0 0 0 32 0 4 2 0 0 0 0 0 0 0 89 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 134 3 0 0 164 3 0 0 9 0 0 10 80 0 0 0 4 0 0 0 9 64 64 128 4 0 128 0 9 64 64 128 4 0 0 1 9 64 64 128 4 0 128 1 9 64 64 128 4 0 0 2 9 128 64 128 5 192 0 0 68 0 128 2 75 0 193 0 92 0 0 1 28 0 1 0 22 0 1 128 70 65 65 2 23 128 193 2 22 64 0 128 75 193 65 2 92 65 0 1 33 128 0 0 22 0 254 127 5 192 0 0 68 0 0 3 70 0 194 0 132 0 0 3 134 64 66 1 156 128 128 0 193 128 2 0 149 192 0 1 92 0 0 1 28 0 1 0 22 128 10 128 68 1 128 3 70 193 194 2 129 129 1 0 196 1 128 2 92 129 128 1 133 65 3 0 134 129 67 3 193 193 3 0 1 2 4 0 156 129 128 1 73 129 1 134 73 129 192 136 134 65 65 2 139 193 68 3 1 194 3 0 65 2 5 0 156 129 0 2 73 129 1 137 73 129 197 138 133 1 6 0 134 65 70 3 193 129 6 0 1 130 6 0 65 130 6 0 156 129 0 2 73 129 129 139 133 1 6 0 134 65 70 3 193 129 6 0 1 130 6 0 65 130 6 0 156 129 0 2 73 129 129 141 134 1 199 2 139 65 71 3 36 2 0 0 4 0 128 2 0 0 128 2 4 0 0 4 0 0 0 2 156 65 128 1 99 1 0 0 227 0 0 0 33 128 0 0 22 128 244 127 30 0 128 0 30 0 0 0 4 8 0 0 0 0 0 0 0 86 105 115 105 98 108 101 0 1 0 1 1 4 6 0 0 0 0 0 0 0 112 97 105 114 115 0 4 12 0 0 0 0 0 0 0 71 101 116 67 104 105 108 100 114 101 110 0 4 5 0 0 0 0 0 0 0 78 97 109 101 0 4 11 0 0 0 0 0 0 0 84 101 120 116 66 117 116 116 111 110 0 4 8 0 0 0 0 0 0 0 68 101 115 116 114 111 121 0 4 9 0 0 0 0 0 0 0 71 101 116 70 105 108 101 115 0 4 17 0 0 0 0 0 0 0 71 101 116 79 83 68 114 105 118 101 76 101 116 116 101 114 0 4 34 0 0 0 0 0 0 0 58 47 83 121 115 116 101 109 47 65 112 112 68 97 116 97 47 66 117 105 108 100 66 114 101 97 107 47 115 97 118 101 115 0 4 9 0 0 0 0 0 0 0 67 114 101 97 116 101 85 73 0 4 5 0 0 0 0 0 0 0 83 105 122 101 0 4 6 0 0 0 0 0 0 0 85 68 105 109 50 0 4 10 0 0 0 0 0 0 0 102 114 111 109 83 99 97 108 101 0 3 0 0 0 0 0 0 240 63 3 154 153 153 153 153 153 201 63 4 11 0 0 0 0 0 0 0 84 101 120 116 83 99 97 108 101 100 0 4 5 0 0 0 0 0 0 0 84 101 120 116 0 4 4 0 0 0 0 0 0 0 115 117 98 0 3 0 0 0 0 0 0 20 192 4 23 0 0 0 0 0 0 0 66 97 99 107 103 114 111 117 110 100 84 114 97 110 115 112 97 114 101 110 99 121 0 3 102 102 102 102 102 102 230 63 4 17 0 0 0 0 0 0 0 66 97 99 107 103 114 111 117 110 100 67 111 108 111 114 51 0 4 7 0 0 0 0 0 0 0 67 111 108 111 114 51 0 4 8 0 0 0 0 0 0 0 102 114 111 109 82 71 66 0 3 0 0 0 0 0 224 111 64 4 11 0 0 0 0 0 0 0 84 101 120 116 67 111 108 111 114 51 0 4 18 0 0 0 0 0 0 0 77 111 117 115 101 66 117 116 116 111 110 49 67 108 105 99 107 0 4 8 0 0 0 0 0 0 0 67 111 110 110 101 99 116 0 1 0 0 0 0 0 0 0 0 0 0 0 154 3 0 0 162 3 0 0 4 0 0 9 30 0 0 0 5 0 0 0 68 0 0 0 75 64 192 0 92 0 0 1 28 0 1 0 22 64 2 128 70 129 64 2 23 192 192 2 22 128 1 128 69 65 1 0 70 129 193 2 129 193 1 0 193 193 1 0 1 194 1 0 92 129 0 2 9 65 1 130 33 128 0 0 22 192 252 127 4 0 128 0 69 64 1 0 70 128 193 0 129 0 2 0 193 0 2 0 1 1 2 0 92 128 0 2 9 64 0 130 4 0 128 1 6 128 64 0 8 0 0 1 30 0 128 0 9 0 0 0 4 6 0 0 0 0 0 0 0 112 97 105 114 115 0 4 12 0 0 0 0 0 0 0 71 101 116 67 104 105 108 100 114 101 110 0 4 5 0 0 0 0 0 0 0 78 97 109 101 0 4 11 0 0 0 0 0 0 0 84 101 120 116 66 117 116 116 111 110 0 4 17 0 0 0 0 0 0 0 66 97 99 107 103 114 111 117 110 100 67 111 108 111 114 51 0 4 7 0 0 0 0 0 0 0 67 111 108 111 114 51 0 4 8 0 0 0 0 0 0 0 102 114 111 109 82 71 66 0 3 0 0 0 0 0 224 111 64 3 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 166 3 0 0 178 3 0 0 9 0 0 6 38 0 0 0 4 0 0 0 69 64 0 0 70 0 192 0 70 128 192 0 9 64 0 128 4 0 0 0 9 0 193 129 4 0 128 0 65 64 1 0 28 64 0 1 4 0 0 1 9 192 65 131 4 0 128 1 9 0 65 131 4 0 0 2 9 0 65 131 4 0 128 2 9 0 65 131 4 0 128 0 65 0 2 0 28 64 0 1 4 0 0 3 28 64 128 0 4 0 128 0 65 64 2 0 28 64 0 1 4 0 128 3 69 128 2 0 70 192 194 0 133 0 3 0 134 192 66 1 196 0 0 4 1 65 3 0 68 1 0 4 156 0 0 2 92 128 0 0 9 64 0 133 30 0 128 0 14 0 0 0 4 14 0 0 0 0 0 0 0 77 111 117 115 101 66 101 104 97 118 105 111 114 0 4 5 0 0 0 0 0 0 0 69 110 117 109 0 4 20 0 0 0 0 0 0 0 76 111 99 107 67 117 114 114 101 110 116 80 111 115 105 116 105 111 110 0 4 17 0 0 0 0 0 0 0 77 111 117 115 101 73 99 111 110 69 110 97 98 108 101 100 0 1 0 4 12 0 0 0 0 0 0 0 99 111 110 102 105 103 32 100 111 110 101 0 4 8 0 0 0 0 0 0 0 86 105 115 105 98 108 101 0 1 1 4 13 0 0 0 0 0 0 0 103 97 109 101 32 118 105 115 105 98 108 101 0 4 13 0 0 0 0 0 0 0 114 101 110 100 101 114 32 115 101 116 117 112 0 4 7 0 0 0 0 0 0 0 67 70 114 97 109 101 0 4 4 0 0 0 0 0 0 0 110 101 119 0 4 8 0 0 0 0 0 0 0 86 101 99 116 111 114 51 0 3 0 0 0 0 0 0 94 64 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 182 3 0 0 189 3 0 0 4 0 0 4 16 0 0 0 4 0 0 0 23 0 64 0 22 0 0 128 30 0 128 0 4 0 0 0 11 64 64 0 129 128 0 0 193 192 0 0 28 128 0 2 8 0 128 0 4 0 0 1 68 0 0 0 28 64 0 1 4 0 128 1 28 64 128 0 30 0 128 0 4 0 0 0 4 1 0 0 0 0 0 0 0 0 4 4 0 0 0 0 0 0 0 115 117 98 0 3 0 0 0 0 0 0 240 63 3 0 0 0 0 0 0 20 192 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 191 3 0 0 194 3 0 0 2 0 0 2 5 0 0 0 4 0 0 0 9 64 64 128 4 0 128 0 9 128 64 128 30 0 128 0 3 0 0 0 4 8 0 0 0 0 0 0 0 86 105 115 105 98 108 101 0 1 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 196 3 0 0 209 3 0 0 14 0 0 2 46 0 0 0 4 0 0 0 9 64 64 128 4 0 128 0 9 128 64 128 4 0 128 1 6 192 64 0 8 0 0 1 5 0 1 0 68 0 128 2 70 192 192 0 28 128 0 1 26 64 0 0 22 0 0 128 1 64 1 0 8 0 0 2 5 0 1 0 68 0 128 3 70 192 192 0 28 128 0 1 26 64 0 0 22 0 0 128 1 64 1 0 8 0 0 3 5 0 1 0 68 0 0 4 70 192 192 0 28 128 0 1 23 128 65 0 22 128 0 128 1 192 1 0 8 0 128 4 22 128 1 128 5 0 1 0 68 0 0 4 70 192 192 0 28 128 0 1 68 0 0 5 14 64 0 0 8 0 128 4 4 0 128 5 68 0 0 6 70 192 192 0 28 64 0 1 4 0 128 6 28 64 128 0 30 0 128 0 8 0 0 0 4 8 0 0 0 0 0 0 0 86 105 115 105 98 108 101 0 1 0 1 1 4 5 0 0 0 0 0 0 0 84 101 120 116 0 4 9 0 0 0 0 0 0 0 116 111 110 117 109 98 101 114 0 3 0 0 0 0 0 128 70 64 0 3 0 0 0 0 0 0 94 64 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 211 3 0 0 217 3 0 0 5 0 0 2 15 0 0 0 4 0 0 0 68 0 128 0 28 64 0 1 4 0 0 1 69 64 0 0 70 0 192 0 70 128 192 0 9 64 0 128 4 0 0 1 9 0 193 129 4 0 128 1 9 128 193 130 4 0 0 2 9 0 193 130 30 0 128 0 7 0 0 0 4 14 0 0 0 0 0 0 0 77 111 117 115 101 66 101 104 97 118 105 111 114 0 4 5 0 0 0 0 0 0 0 69 110 117 109 0 4 20 0 0 0 0 0 0 0 76 111 99 107 67 117 114 114 101 110 116 80 111 115 105 116 105 111 110 0 4 17 0 0 0 0 0 0 0 77 111 117 115 101 73 99 111 110 69 110 97 98 108 101 100 0 1 0 4 8 0 0 0 0 0 0 0 86 105 115 105 98 108 101 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 219 3 0 0 227 3 0 0 5 0 0 2 19 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 4 0 128 0 26 0 0 0 22 128 0 128 4 0 128 0 11 64 64 0 28 64 0 1 4 0 0 1 11 64 64 0 28 64 0 1 4 0 128 1 11 64 64 0 28 64 0 1 4 0 0 2 11 64 64 0 28 64 0 1 30 0 128 0 2 0 0 0 4 23 0 0 0 0 0 0 0 98 117 105 108 100 98 114 101 97 107 32 100 105 115 99 111 110 110 101 99 116 115 0 4 11 0 0 0 0 0 0 0 68 105 115 99 111 110 110 101 99 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 