LEF            PaleNoobs                       e61a4f7f2f8337fd68c95374360256efa33706c8bf2abfe97b4871fb34c0f6f5LuaQ         @                 A@  @  �           print        Hello, world!                            