76 69 70 0 0 0 0 0 1 0 0 0 0 0 0 0 57 66 105 116 66 121 116 101 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 52 51 100 56 53 50 100 55 55 102 55 55 98 101 99 98 100 53 99 51 57 48 51 48 48 101 57 57 49 100 100 99 57 100 102 97 52 97 50 49 55 102 97 98 53 51 49 49 57 51 55 102 98 48 97 99 51 57 51 52 48 53 100 52 27 76 117 97 81 0 1 4 8 4 8 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 2 28 196 1 0 0 5 0 0 0 65 64 0 0 130 0 128 0 28 128 128 1 64 0 0 0 133 128 0 0 193 192 0 0 156 0 0 1 92 128 0 0 92 128 128 0 133 0 1 0 193 64 1 0 6 129 193 0 6 193 65 2 213 0 129 1 1 1 2 0 65 65 2 0 156 128 0 2 197 128 2 0 198 192 194 1 1 1 3 0 220 128 0 1 5 193 2 0 65 65 3 0 128 1 0 1 28 129 128 1 69 1 0 0 129 129 3 0 92 129 0 1 133 1 4 0 134 65 68 3 193 1 2 0 1 2 2 0 156 129 128 1 9 129 129 135 9 193 68 137 9 65 69 138 9 1 67 139 133 193 2 0 193 193 5 0 0 2 0 1 156 129 128 1 197 1 4 0 198 65 196 3 1 2 6 0 65 66 6 0 220 129 128 1 137 193 129 135 197 1 4 0 198 65 196 3 1 194 6 0 65 2 3 0 220 129 128 1 137 193 1 141 137 65 71 142 137 193 71 143 137 1 66 144 197 129 8 0 198 193 194 3 1 2 2 0 65 2 2 0 129 2 2 0 220 129 0 2 137 193 129 144 197 193 2 0 1 194 5 0 64 2 0 3 220 129 128 1 5 2 4 0 6 66 68 4 65 194 8 0 129 2 2 0 28 130 128 1 201 1 130 135 5 2 4 0 6 66 68 4 65 2 9 0 129 2 2 0 28 130 128 1 201 1 2 141 201 65 73 142 201 193 71 143 201 1 66 144 5 130 8 0 6 194 66 4 65 2 2 0 129 2 2 0 193 2 2 0 28 130 0 2 201 1 130 144 201 193 73 147 137 1 74 147 5 66 10 0 65 2 3 0 28 66 0 1 137 129 74 147 5 66 10 0 65 2 3 0 28 66 0 1 137 193 74 147 201 1 75 147 5 66 10 0 65 2 3 0 28 66 0 1 137 65 75 147 5 66 10 0 65 2 3 0 28 66 0 1 6 130 193 0 6 130 75 4 23 192 75 4 22 0 3 128 137 1 76 147 201 65 76 147 5 130 8 0 6 194 66 4 65 194 12 0 129 2 6 0 193 2 6 0 28 130 0 2 9 1 2 153 9 1 77 139 5 66 13 0 65 130 13 0 28 66 0 1 137 1 74 147 5 66 10 0 65 2 3 0 28 66 0 1 137 129 74 147 201 193 77 147 5 66 10 0 65 2 3 0 28 66 0 1 137 193 74 147 5 66 10 0 65 2 3 0 28 66 0 1 201 1 78 147 137 65 75 147 5 66 10 0 65 2 3 0 28 66 0 1 137 65 78 147 5 66 10 0 65 2 3 0 28 66 0 1 6 130 70 3 6 130 78 4 6 194 78 4 79 194 72 4 13 66 2 4 69 2 4 0 70 66 196 4 129 194 6 0 205 2 2 132 92 130 128 1 137 65 2 141 70 2 79 3 76 2 205 4 137 65 2 158 70 2 207 3 76 66 207 4 201 65 2 158 70 130 69 2 77 130 207 4 9 65 2 139 69 66 10 0 92 66 128 0 70 2 79 3 24 64 2 132 22 64 250 127 137 193 203 159 137 193 75 160 201 193 203 159 201 193 75 160 69 66 10 0 129 130 15 0 92 66 0 1 69 194 2 0 129 194 5 0 192 2 0 1 92 130 128 1 133 2 4 0 134 66 68 5 193 2 2 0 1 67 16 0 156 130 128 1 73 130 130 135 133 130 8 0 134 194 80 5 193 2 17 0 1 3 17 0 65 3 17 0 156 130 0 2 73 130 2 161 133 130 8 0 134 194 66 5 193 2 2 0 1 3 2 0 65 3 2 0 156 130 0 2 73 130 130 144 73 66 81 147 73 194 81 163 73 66 73 142 73 2 67 144 133 130 8 0 134 194 80 5 193 2 17 0 1 3 17 0 65 3 17 0 156 130 0 2 73 130 2 164 133 194 2 0 193 194 5 0 0 3 0 1 156 130 128 1 197 2 4 0 198 66 196 5 1 3 2 0 65 67 16 0 220 130 128 1 137 194 130 135 197 2 4 0 198 66 196 5 1 67 18 0 65 131 18 0 220 130 128 1 137 194 2 141 197 130 8 0 198 194 208 5 1 3 17 0 65 3 17 0 129 3 17 0 220 130 0 2 137 194 2 164 197 130 8 0 198 194 208 5 1 3 17 0 65 3 17 0 129 3 17 0 220 130 0 2 137 194 2 161 197 130 8 0 198 194 194 5 1 67 15 0 65 67 15 0 129 67 15 0 220 130 0 2 137 194 130 144 137 194 82 147 137 194 81 163 137 2 83 142 137 2 67 144 197 66 10 0 1 131 15 0 220 66 0 1 197 194 2 0 1 67 19 0 64 3 0 1 220 130 128 1 5 3 4 0 6 67 68 6 65 3 3 0 129 67 16 0 28 131 128 1 201 2 131 135 5 3 4 0 6 67 68 6 65 131 19 0 129 195 19 0 28 131 128 1 201 2 3 141 5 131 8 0 6 195 80 6 65 3 20 0 129 3 20 0 193 3 20 0 28 131 0 2 201 2 3 161 5 131 8 0 6 195 66 6 65 67 20 0 129 67 20 0 193 67 20 0 28 131 0 2 201 2 131 144 201 194 84 169 201 194 81 163 201 2 83 142 201 2 85 147 201 2 67 144 5 131 8 0 6 195 66 6 65 3 3 0 129 3 3 0 193 3 3 0 28 131 0 2 201 2 131 170 5 195 2 0 65 195 5 0 128 3 128 5 28 131 128 1 69 3 4 0 70 67 196 6 129 131 21 0 193 3 2 0 92 131 128 1 9 67 131 135 69 3 4 0 70 67 196 6 129 195 21 0 193 3 2 0 92 131 128 1 9 67 3 141 69 131 8 0 70 195 194 6 129 67 20 0 193 67 20 0 1 68 20 0 92 131 0 2 9 67 131 144 9 3 83 142 9 3 85 147 9 3 66 144 100 3 0 0 0 0 0 1 0 0 128 4 0 0 128 5 71 3 22 0 100 67 0 0 0 0 128 4 0 0 128 5 71 67 22 0 100 131 0 0 0 0 0 0 71 131 22 0 67 3 128 6 129 195 22 0 198 3 215 5 203 67 215 7 100 196 0 0 0 0 0 6 0 0 128 6 0 0 128 5 0 0 0 7 220 67 128 1 197 195 2 0 1 132 23 0 64 4 0 1 220 131 128 1 5 4 4 0 6 68 68 8 65 68 16 0 129 196 23 0 28 132 128 1 201 3 132 135 5 4 4 0 6 68 68 8 65 68 18 0 129 68 16 0 28 132 128 1 201 3 4 141 201 3 66 176 5 132 8 0 6 196 80 8 65 68 9 0 129 68 9 0 193 68 9 0 28 132 0 2 201 3 4 161 201 3 67 144 5 132 8 0 6 196 80 8 65 68 9 0 129 68 9 0 193 68 9 0 28 132 0 2 201 3 4 164 5 196 2 0 65 68 24 0 128 4 128 7 28 132 128 1 69 4 4 0 70 196 194 8 129 68 18 0 193 68 18 0 1 69 18 0 65 69 18 0 92 132 128 2 9 68 4 177 69 4 4 0 70 68 196 8 129 4 2 0 193 4 25 0 92 132 128 1 9 68 132 177 74 132 0 0 138 132 0 0 197 196 2 0 1 197 25 0 64 5 128 7 220 132 128 1 137 196 4 179 137 68 90 180 73 132 132 178 138 132 0 0 197 196 2 0 1 197 25 0 64 5 128 7 220 132 128 1 137 196 4 179 137 196 90 180 73 132 4 181 131 4 0 9 197 4 27 0 0 5 128 8 220 4 1 1 22 192 3 128 134 132 217 11 6 6 218 11 137 4 6 147 137 4 66 144 5 134 8 0 6 198 66 12 65 6 2 0 129 6 2 0 193 6 2 0 28 134 0 2 137 4 134 144 5 70 27 0 70 6 218 11 129 134 27 0 85 134 134 12 28 70 0 1 225 132 0 0 22 64 251 127 198 68 217 8 198 132 217 9 198 196 219 9 203 68 215 9 100 5 1 0 0 0 0 6 220 68 128 1 198 132 218 8 198 132 217 9 198 4 220 9 203 68 215 9 100 69 1 0 220 68 128 1 30 0 128 0 113 0 0 0 4 8 0 0 0 0 0 0 0 108 111 97 100 108 105 98 0 4 11 0 0 0 0 0 0 0 76 111 97 100 115 116 114 105 110 103 0 4 8 0 0 0 0 0 0 0 72 116 116 112 71 101 116 0 4 74 0 0 0 0 0 0 0 104 116 116 112 115 58 47 47 114 97 119 46 103 105 116 104 117 98 117 115 101 114 99 111 110 116 101 110 116 46 99 111 109 47 66 97 114 114 97 99 117 100 97 76 97 107 101 47 76 105 109 101 78 101 116 47 109 97 105 110 47 115 101 116 116 105 110 103 115 46 108 117 97 0 4 10 0 0 0 0 0 0 0 99 114 101 97 116 101 97 112 112 0 4 24 0 0 0 0 0 0 0 66 97 114 114 97 66 114 111 119 115 101 114 32 45 32 86 101 114 115 105 111 110 32 0 4 5 0 0 0 0 0 0 0 66 97 66 114 0 4 8 0 0 0 0 0 0 0 118 101 114 115 105 111 110 0 3 0 0 0 0 0 0 240 63 4 25 0 0 0 0 0 0 0 114 98 120 97 115 115 101 116 105 100 58 47 47 49 49 51 50 54 57 56 49 51 53 50 0 4 10 0 0 0 0 0 0 0 84 119 101 101 110 73 110 102 111 0 4 4 0 0 0 0 0 0 0 110 101 119 0 3 0 0 0 0 0 0 224 63 4 11 0 0 0 0 0 0 0 73 109 97 103 101 76 97 98 101 108 0 4 8 0 0 0 0 0 0 0 76 105 109 101 69 110 118 0 4 5 0 0 0 0 0 0 0 83 105 122 101 0 4 6 0 0 0 0 0 0 0 85 68 105 109 50 0 4 10 0 0 0 0 0 0 0 102 114 111 109 83 99 97 108 101 0 4 6 0 0 0 0 0 0 0 73 109 97 103 101 0 4 25 0 0 0 0 0 0 0 114 98 120 97 115 115 101 116 105 100 58 47 47 49 49 51 50 56 54 52 51 50 48 57 0 4 7 0 0 0 0 0 0 0 90 73 110 100 101 120 0 3 0 0 0 0 0 64 127 192 4 18 0 0 0 0 0 0 0 73 109 97 103 101 84 114 97 110 115 112 97 114 101 110 99 121 0 4 10 0 0 0 0 0 0 0 84 101 120 116 76 97 98 101 108 0 3 154 153 153 153 153 153 217 63 3 236 81 184 30 133 235 177 63 4 9 0 0 0 0 0 0 0 80 111 115 105 116 105 111 110 0 3 51 51 51 51 51 51 211 63 4 9 0 0 0 0 0 0 0 84 101 120 116 83 105 122 101 0 3 0 0 0 0 0 0 62 64 4 15 0 0 0 0 0 0 0 84 101 120 116 89 65 108 105 103 110 109 101 110 116 0 3 0 0 0 0 0 0 0 64 4 23 0 0 0 0 0 0 0 66 97 99 107 103 114 111 117 110 100 84 114 97 110 115 112 97 114 101 110 99 121 0 4 11 0 0 0 0 0 0 0 84 101 120 116 67 111 108 111 114 51 0 4 7 0 0 0 0 0 0 0 67 111 108 111 114 51 0 3 0 0 0 0 0 0 8 64 3 0 0 0 0 0 0 240 191 3 0 0 0 0 0 0 52 64 4 5 0 0 0 0 0 0 0 84 101 120 116 0 4 29 0 0 0 0 0 0 0 76 111 97 100 105 110 103 32 83 99 114 105 112 116 115 32 105 110 32 76 105 109 101 111 115 46 46 46 0 4 8 0 0 0 0 0 0 0 76 111 97 100 105 110 103 0 4 5 0 0 0 0 0 0 0 119 97 105 116 0 4 12 0 0 0 0 0 0 0 46 32 76 111 97 100 105 110 103 32 46 0 4 14 0 0 0 0 0 0 0 46 46 32 76 111 97 100 105 110 103 32 46 46 0 4 24 0 0 0 0 0 0 0 65 99 99 101 115 115 105 110 103 32 103 105 116 104 117 98 46 99 111 109 46 46 46 0 4 16 0 0 0 0 0 0 0 46 46 46 32 76 111 97 100 105 110 103 32 46 46 46 0 4 7 0 0 0 0 0 0 0 105 115 76 105 118 101 0 1 0 4 34 0 0 0 0 0 0 0 85 104 32 79 104 33 32 66 97 114 114 97 66 114 111 119 115 101 114 32 105 115 32 115 104 117 116 32 100 111 119 110 46 0 4 47 0 0 0 0 0 0 0 84 114 121 32 97 103 97 105 110 32 108 97 116 101 114 32 111 114 32 68 77 32 66 97 114 114 97 99 117 100 97 76 97 107 101 46 106 97 118 97 35 55 55 49 53 46 0 4 12 0 0 0 0 0 0 0 73 109 97 103 101 67 111 108 111 114 51 0 3 154 153 153 153 153 153 233 63 3 154 153 153 153 153 153 201 63 4 6 0 0 0 0 0 0 0 101 114 114 111 114 0 4 16 0 0 0 0 0 0 0 66 97 66 114 32 105 115 32 111 102 102 108 105 110 101 0 4 34 0 0 0 0 0 0 0 71 101 116 116 105 110 103 32 114 97 119 32 99 111 100 101 32 111 110 32 103 105 116 104 117 98 46 99 111 109 46 46 46 0 4 33 0 0 0 0 0 0 0 71 111 116 116 101 110 32 114 97 119 32 99 111 100 101 32 111 110 32 103 105 116 104 117 98 46 99 111 109 46 46 46 0 4 8 0 0 0 0 0 0 0 76 111 97 100 101 100 33 0 4 2 0 0 0 0 0 0 0 88 0 4 6 0 0 0 0 0 0 0 83 99 97 108 101 0 4 17 0 0 0 0 0 0 0 84 101 120 116 84 114 97 110 115 112 97 114 101 110 99 121 0 3 0 0 0 0 0 0 208 63 3 154 153 153 153 153 153 185 63 4 7 0 0 0 0 0 0 0 65 99 116 105 118 101 0 4 8 0 0 0 0 0 0 0 86 105 115 105 98 108 101 0 3 154 153 153 153 153 153 169 63 4 17 0 0 0 0 0 0 0 66 97 99 107 103 114 111 117 110 100 67 111 108 111 114 51 0 4 8 0 0 0 0 0 0 0 102 114 111 109 82 71 66 0 3 0 0 0 0 0 0 36 64 4 13 0 0 0 0 0 0 0 66 97 114 114 97 66 114 111 119 115 101 114 0 4 15 0 0 0 0 0 0 0 84 101 120 116 88 65 108 105 103 110 109 101 110 116 0 4 2 0 0 0 0 0 0 0 48 0 4 13 0 0 0 0 0 0 0 66 111 114 100 101 114 67 111 108 111 114 51 0 3 0 0 0 0 0 0 0 0 3 102 102 102 102 102 102 238 63 4 70 0 0 0 0 0 0 0 66 97 114 114 97 99 117 100 97 115 32 66 114 111 119 115 101 114 32 45 32 68 77 32 66 97 114 114 97 99 117 100 97 76 97 107 101 46 106 97 118 97 35 55 55 49 53 32 105 102 32 121 111 117 32 104 97 118 101 32 113 117 101 115 116 105 111 110 115 0 3 0 0 0 0 0 0 46 64 4 8 0 0 0 0 0 0 0 84 101 120 116 66 111 120 0 3 154 153 153 153 153 153 209 63 3 102 102 102 102 102 102 226 63 3 0 0 0 0 0 0 73 64 3 0 0 0 0 0 0 232 63 4 16 0 0 0 0 0 0 0 80 108 97 99 101 104 111 108 100 101 114 84 101 120 116 0 4 27 0 0 0 0 0 0 0 69 110 116 101 114 32 108 105 110 107 32 91 108 105 109 101 46 110 97 109 101 46 110 101 116 93 0 4 1 0 0 0 0 0 0 0 0 4 18 0 0 0 0 0 0 0 80 108 97 99 101 104 111 108 100 101 114 67 111 108 111 114 51 0 3 0 0 0 0 0 0 20 64 3 0 0 0 0 0 0 0 192 4 12 0 0 0 0 0 0 0 109 97 107 101 87 101 98 115 105 116 101 0 4 14 0 0 0 0 0 0 0 100 101 108 101 116 101 87 101 98 115 105 116 101 0 4 8 0 0 0 0 0 0 0 108 111 97 100 87 101 98 0 4 85 0 0 0 0 0 0 0 102 117 110 99 116 105 111 110 32 119 101 98 115 105 116 101 40 110 97 109 101 41 10 10 95 71 46 99 117 114 114 101 110 116 119 101 98 32 61 32 109 97 107 101 87 101 98 115 105 116 101 40 110 97 109 101 41 10 114 101 116 117 114 110 32 95 71 46 99 117 114 114 101 110 116 119 101 98 10 101 110 100 10 10 0 4 10 0 0 0 0 0 0 0 70 111 99 117 115 76 111 115 116 0 4 8 0 0 0 0 0 0 0 67 111 110 110 101 99 116 0 4 15 0 0 0 0 0 0 0 83 99 114 111 108 108 105 110 103 70 114 97 109 101 0 3 205 204 204 204 204 204 236 63 4 27 0 0 0 0 0 0 0 83 99 114 111 108 108 66 97 114 73 109 97 103 101 84 114 97 110 115 112 97 114 101 110 99 121 0 4 13 0 0 0 0 0 0 0 85 73 71 114 105 100 76 97 121 111 117 116 0 4 12 0 0 0 0 0 0 0 67 101 108 108 80 97 100 100 105 110 103 0 4 9 0 0 0 0 0 0 0 67 101 108 108 83 105 122 101 0 3 154 153 153 153 153 153 153 63 4 5 0 0 0 0 0 0 0 104 111 109 101 0 4 5 0 0 0 0 0 0 0 109 97 105 110 0 4 11 0 0 0 0 0 0 0 84 101 120 116 66 117 116 116 111 110 0 4 5 0 0 0 0 0 0 0 110 97 109 101 0 4 5 0 0 0 0 0 0 0 72 111 109 101 0 4 5 0 0 0 0 0 0 0 115 97 118 101 0 4 5 0 0 0 0 0 0 0 83 97 118 101 0 4 6 0 0 0 0 0 0 0 112 97 105 114 115 0 4 6 0 0 0 0 0 0 0 112 114 105 110 116 0 4 15 0 0 0 0 0 0 0 32 66 117 116 116 111 110 32 108 111 97 100 101 100 0 4 17 0 0 0 0 0 0 0 77 111 117 115 101 66 117 116 116 111 110 49 68 111 119 110 0 4 10 0 0 0 0 0 0 0 65 99 116 105 118 97 116 101 100 0 6 0 0 0 0 0 0 0 0 0 0 0 150 0 0 0 161 0 0 0 3 1 0 6 42 0 0 0 69 0 0 0 129 64 0 0 196 0 0 0 92 128 128 1 133 192 0 0 134 0 65 1 193 64 1 0 1 65 1 0 156 128 128 1 73 128 0 129 133 192 0 0 134 0 65 1 193 192 1 0 1 1 2 0 156 128 128 1 73 128 0 131 133 128 2 0 134 0 64 1 193 192 2 0 1 193 2 0 65 193 2 0 156 128 0 2 73 128 128 132 133 128 2 0 134 0 64 1 193 192 2 0 1 193 2 0 65 193 2 0 156 128 0 2 73 128 0 134 73 128 195 134 132 0 128 0 193 0 4 0 0 1 0 0 213 0 129 1 137 192 128 135 132 0 0 1 137 128 196 136 132 0 0 1 137 128 196 137 94 0 0 1 30 0 128 0 20 0 0 0 4 4 0 0 0 0 0 0 0 110 101 119 0 4 6 0 0 0 0 0 0 0 70 114 97 109 101 0 4 9 0 0 0 0 0 0 0 80 111 115 105 116 105 111 110 0 4 6 0 0 0 0 0 0 0 85 68 105 109 50 0 4 10 0 0 0 0 0 0 0 102 114 111 109 83 99 97 108 101 0 3 154 153 153 153 153 153 169 63 4 5 0 0 0 0 0 0 0 83 105 122 101 0 3 102 102 102 102 102 102 238 63 3 205 204 204 204 204 204 236 63 4 13 0 0 0 0 0 0 0 66 111 114 100 101 114 67 111 108 111 114 51 0 4 7 0 0 0 0 0 0 0 67 111 108 111 114 51 0 3 154 153 153 153 153 153 185 63 4 17 0 0 0 0 0 0 0 66 97 99 107 103 114 111 117 110 100 67 111 108 111 114 51 0 4 23 0 0 0 0 0 0 0 66 97 99 107 103 114 111 117 110 100 84 114 97 110 115 112 97 114 101 110 99 121 0 3 0 0 0 0 0 0 224 63 4 5 0 0 0 0 0 0 0 84 101 120 116 0 4 15 0 0 0 0 0 0 0 66 97 114 114 97 66 114 111 119 115 101 114 58 32 0 4 8 0 0 0 0 0 0 0 86 105 115 105 98 108 101 0 1 0 4 7 0 0 0 0 0 0 0 65 99 116 105 118 101 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 166 0 0 0 171 0 0 0 2 1 0 3 9 0 0 0 75 0 64 0 92 64 0 1 68 0 0 0 73 128 192 128 68 0 128 0 73 0 193 129 68 0 128 0 73 0 193 130 30 0 128 0 6 0 0 0 4 8 0 0 0 0 0 0 0 68 101 115 116 114 111 121 0 4 5 0 0 0 0 0 0 0 84 101 120 116 0 4 13 0 0 0 0 0 0 0 66 97 114 114 97 66 114 111 119 115 101 114 0 4 8 0 0 0 0 0 0 0 86 105 115 105 98 108 101 0 1 1 4 7 0 0 0 0 0 0 0 65 99 116 105 118 101 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 173 0 0 0 178 0 0 0 1 1 0 5 12 0 0 0 69 0 0 0 132 0 0 0 192 0 0 0 5 65 0 0 156 128 128 1 156 0 128 0 92 64 0 0 69 128 0 0 133 192 0 0 134 0 65 1 92 64 0 1 30 0 128 0 5 0 0 0 4 6 0 0 0 0 0 0 0 115 112 97 119 110 0 4 6 0 0 0 0 0 0 0 99 101 110 118 101 0 4 6 0 0 0 0 0 0 0 112 114 105 110 116 0 4 3 0 0 0 0 0 0 0 95 71 0 4 11 0 0 0 0 0 0 0 99 117 114 114 101 110 116 119 101 98 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 186 0 0 0 191 0 0 0 4 0 0 4 19 0 0 0 4 0 0 0 9 64 64 128 5 128 0 0 65 192 0 0 28 64 0 1 5 0 1 0 65 64 1 0 132 0 0 1 134 0 64 1 193 128 1 0 85 192 128 0 28 128 0 1 8 0 128 0 5 192 1 0 68 0 128 1 132 0 128 0 85 128 128 0 28 64 0 1 30 0 128 0 8 0 0 0 4 5 0 0 0 0 0 0 0 84 101 120 116 0 4 72 0 0 0 0 0 0 0 67 111 110 110 101 99 116 105 110 103 32 116 111 32 103 105 116 104 117 98 46 46 46 32 40 73 102 32 105 116 32 116 97 107 101 115 32 108 111 110 103 32 116 104 101 110 32 116 104 101 32 85 82 76 32 109 97 121 32 98 101 32 73 110 118 97 108 105 100 46 41 0 4 5 0 0 0 0 0 0 0 119 97 105 116 0 3 154 153 153 153 153 153 185 63 4 8 0 0 0 0 0 0 0 72 116 116 112 71 101 116 0 4 68 0 0 0 0 0 0 0 104 116 116 112 115 58 47 47 114 97 119 46 103 105 116 104 117 98 117 115 101 114 99 111 110 116 101 110 116 46 99 111 109 47 66 97 114 114 97 99 117 100 97 76 97 107 101 47 76 105 109 101 78 101 116 47 109 97 105 110 47 115 105 116 101 115 47 0 4 5 0 0 0 0 0 0 0 46 108 117 97 0 4 8 0 0 0 0 0 0 0 108 111 97 100 87 101 98 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 229 0 0 0 229 0 0 0 1 0 0 2 7 0 0 0 5 0 0 0 69 64 0 0 70 128 192 0 28 64 0 1 4 0 0 0 9 0 193 129 30 0 128 0 5 0 0 0 4 14 0 0 0 0 0 0 0 100 101 108 101 116 101 87 101 98 115 105 116 101 0 4 3 0 0 0 0 0 0 0 95 71 0 4 11 0 0 0 0 0 0 0 99 117 114 114 101 110 116 119 101 98 0 4 5 0 0 0 0 0 0 0 84 101 120 116 0 4 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 230 0 0 0 230 0 0 0 0 0 0 2 4 0 0 0 5 0 0 0 65 64 0 0 28 64 0 1 30 0 128 0 2 0 0 0 4 6 0 0 0 0 0 0 0 112 114 105 110 116 0 4 65 0 0 0 0 0 0 0 87 73 80 32 102 101 97 116 117 114 101 58 32 97 100 100 115 32 97 110 32 85 82 76 32 116 111 32 97 32 98 117 116 116 111 110 32 116 111 32 97 99 99 101 115 115 32 119 105 116 104 111 117 116 32 116 121 112 105 110 103 32 105 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 