76 69 70 0 0 0 0 0 1 0 0 0 0 0 0 0 57 66 105 116 66 121 116 101 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 52 49 54 102 51 102 55 102 102 56 50 50 54 51 53 48 49 48 101 101 98 98 100 57 53 100 52 51 50 98 48 55 101 101 101 54 50 99 51 54 55 52 101 98 51 56 56 55 99 99 50 51 48 56 54 51 54 99 48 57 53 97 48 50 27 76 117 97 81 0 1 4 8 4 8 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 2 3 13 0 0 0 5 0 0 0 6 64 64 0 65 128 0 0 28 64 0 1 5 192 0 0 69 0 1 0 129 64 1 0 92 128 0 1 70 128 193 0 133 192 1 0 92 0 0 1 28 64 0 0 30 0 128 0 8 0 0 0 4 5 0 0 0 0 0 0 0 76 105 109 101 0 4 13 0 0 0 0 0 0 0 67 114 101 97 116 101 87 105 110 100 111 119 0 4 7 0 0 0 0 0 0 0 104 101 108 108 111 33 0 4 4 0 0 0 0 0 0 0 108 111 103 0 4 8 0 0 0 0 0 0 0 108 111 97 100 108 105 98 0 4 11 0 0 0 0 0 0 0 68 82 77 77 97 110 97 103 101 114 0 4 8 0 0 0 0 0 0 0 79 119 110 115 65 112 112 0 4 7 0 0 0 0 0 0 0 115 99 114 105 112 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 