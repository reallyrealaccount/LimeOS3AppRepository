76 69 70 0 0 0 0 0 1 0 0 0 0 0 0 0 57 66 105 116 66 121 116 101 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 57 55 54 102 52 102 97 102 53 53 56 53 57 97 98 56 49 52 57 49 51 52 98 50 97 99 49 55 99 102 53 53 52 98 55 51 48 55 49 49 51 53 55 57 98 50 99 52 56 97 49 97 99 102 52 51 97 97 99 98 57 54 102 98 27 76 117 97 81 0 1 4 8 4 8 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 2 3 11 0 0 0 5 0 0 0 65 64 0 0 28 128 0 1 69 128 0 0 129 192 0 0 92 128 0 1 133 0 1 0 156 0 128 0 28 128 0 0 28 64 128 0 30 0 128 0 5 0 0 0 4 8 0 0 0 0 0 0 0 108 111 97 100 108 105 98 0 4 11 0 0 0 0 0 0 0 76 111 97 100 115 116 114 105 110 103 0 4 8 0 0 0 0 0 0 0 72 116 116 112 71 101 116 0 4 81 0 0 0 0 0 0 0 104 116 116 112 115 58 47 47 114 97 119 46 103 105 116 104 117 98 117 115 101 114 99 111 110 116 101 110 116 46 99 111 109 47 66 105 103 109 97 110 99 111 122 109 111 47 108 105 109 101 111 115 45 103 97 109 101 45 115 116 117 100 105 111 47 109 97 105 110 47 115 99 114 105 112 116 46 108 117 97 0 4 8 0 0 0 0 0 0 0 103 101 116 102 101 110 118 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 