LEF            ruben070hallo                   3dc6ca3394177c56fbd794eca782f1c1595b91acd44216b5c74921a4761aa17dLuaQ         @           .     A@  ��  ��E�  �  �@A \��I�A��@ � B��BI� �I Å�� ��@�� � A �� ���I����� ��@�� � A� �� ���I����@ ��@�� � A �� I� �I�ƌI ǍI�ǎI�Ï��  �     ���ŀ �@�� A� �� �� ܀�����ŀ ���� A� �� �� ܀������@ ���� A	 �� ܀ ������  A	 @  ܀�� �@A� �� �� � ��� ��� �@A�	 �� �� � ��� ��A �@A� �	 �� � � ��� ʓA B�B� ��@ʍɀJ�ɀǕA �@A� �� � � � ��  A �  ��	�˖E� F����	 ��	 �	 A�	 \��	A��	�ƅF�KK��     \A�FALK��A     \A�F�LK��  \A�E�  � �  \��I�̖�� ��@��	 �	 A�	 ��	 ���I����� ��@��	 � A� �� ���I���I�ƅ����L$�    ��A��A��L$   ��A���  �    ���Ł ���� A� �� �� ܁�������ƅ��K��dB    �A��AL��d�    �A���   @  ܁��͖� �@A�	 ��	 ��	 �	 ������ �@A� �� �� � �����Ɂƅ��L��   �B�B�L�   �B��  A �  ��	B͖E� F����	 ��	 �	 A�	 \��	B��E� F���� �� � A� \��	B��	�ƅF�KK��B    \B�FBLK��    \B�E�  �B	 �  \���� ��@��	 � A� �� ���I����� ��@�� � A� �� ���I����B ��@�� 	 A� �� I���I�Ó�B �B��BI��I�͍I�ƌIΕIBN�IN��B ��@�� � A �� I�� � ;   
       createapp                rbxassetid://9397029482        new 
       TextLabel        Parent        Text        PhotoLime v1        Font        Enum        Ubuntu        ZIndex        @	       Position        UDim2         {�G�z�?       Size ffffff�?�Q���?       TextColor3        Color3 333333�?�������?      �?       BackgroundTransparency       �?	       TextSize       4@       ClipsDescendants        TextXAlignment        Frame 
       fromScale �������?       BackgroundColor3 {�G�z�?       TextButton �������?       BorderSizePixel ������@      D@       Page 1        TextScaled        ImageButton        Image +       http://www.roblox.com/asset/?id=8425069718        MouseEnter        Connect        MouseLeave        MouseButton1Click +       http://www.roblox.com/asset/?id=8345858114 +       http://www.roblox.com/asset/?id=8450601351 +       http://www.roblox.com/asset/?id=6075395846 333333�?      6@        More Soon!        Active            &   )           E@  F�� ��  ��  �  A�  \��	@ �   	@A� �           Size        UDim2        new ��Q��?       ZIndex        @       '   '   '   '   '   '   '   '   '   (   (   )                 Image1         +   .           E@  F�� ��  ��  �  A�  \��	@ �   	@A� �           Size        UDim2        new �������?       ZIndex       �?       ,   ,   ,   ,   ,   ,   ,   ,   ,   -   -   .                 Image1         0   2            @@ @@ @@ �@ �@ 	@A� �           script        Parent        HomeScreen        Background        Image +       http://www.roblox.com/asset/?id=8425069718        1   1   1   1   1   1   1   2                   :   =           E@  F�� ��  ��  �  A�  \��	@ �   	@A� �           Size        UDim2        new ��Q��?       ZIndex        @       ;   ;   ;   ;   ;   ;   ;   ;   ;   <   <   =                 Image2         ?   B           E@  F�� ��  ��  �  A�  \��	@ �   	@A� �           Size        UDim2        new �������?       ZIndex       �?       @   @   @   @   @   @   @   @   @   A   A   B                 Image2         I   L           E@  F�� ��  ��  �  A�  \��	@ �   	@A� �           Size        UDim2        new ��Q��?       ZIndex        @       J   J   J   J   J   J   J   J   J   K   K   L                 Image3         N   Q           E@  F�� ��  ��  �  A�  \��	@ �   	@A� �           Size        UDim2        new �������?       ZIndex       �?       O   O   O   O   O   O   O   O   O   P   P   Q                 Image3         Z   ]           E@  F�� ��  ��  �  A�  \��	@ �   	@A� �           Size        UDim2        new ��Q��?       ZIndex        @       [   [   [   [   [   [   [   [   [   \   \   ]                 Image4         _   b           E@  F�� ��  ��  �  A�  \��	@ �   	@A� �           Size        UDim2        new �������?       ZIndex       �?       `   `   `   `   `   `   `   `   `   a   a   b                 Image4         k   n           E@  F�� ��  ��  �  A�  \��	@ �   	@A� �           Size        UDim2        new ��Q��?       ZIndex        @       l   l   l   l   l   l   l   l   l   m   m   n                 Image5         p   s           E@  F�� ��  ��  �  A�  \��	@ �   	@A� �           Size        UDim2        new �������?       ZIndex       �?       q   q   q   q   q   q   q   q   q   r   r   s                 Image5 .                                            	   	   	   	   	   	   	   	   
   
   
   
   
   
   
   
                                                                                                                                                                                                                                                   !   !   !   !   "   #   #   #   #   #   #   #   #   $   &   &   )   )   &   +   +   .   .   +   0   0   2   0   4   4   4   4   5   6   6   6   6   6   6   6   6   7   7   7   7   7   7   7   7   8   :   :   =   =   :   ?   ?   B   B   ?   D   D   D   D   F   F   F   F   F   F   F   F   G   I   I   L   L   I   N   N   Q   Q   N   T   T   T   T   U   V   V   V   V   V   V   V   V   W   W   W   W   W   W   W   W   X   Z   Z   ]   ]   Z   _   _   b   b   _   e   e   e   e   f   g   g   g   g   g   g   g   g   h   h   h   h   h   h   h   h   i   k   k   n   n   k   p   p   s   s   p   u   u   u   u   v   v   v   v   v   v   v   v   w   w   w   w   w   w   w   w   x   x   x   x   x   x   x   y   z   z   z   z   {   |   }   ~      �   �   �   �   �   �   �   �   
          app    -         AppName    -         bar -   -         HomeButton H   -         Image1 r   -         Image2 �   -         Image3 �   -         Image4 �   -         Image5 �   -         HomeButton2   -      