76 69 70 0 0 0 0 0 1 0 0 0 0 0 0 0 114 117 98 101 110 48 55 48 104 97 108 108 111 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 54 57 99 99 51 52 53 52 52 101 55 101 56 97 57 97 57 97 57 101 52 54 51 50 50 99 102 57 53 102 100 51 102 51 98 100 49 50 49 48 52 100 55 98 51 57 99 56 102 56 99 55 56 101 57 102 52 99 99 53 56 52 50 51 27 76 117 97 81 0 1 4 8 4 8 0 2 0 0 0 0 0 0 0 64 0 0 0 0 0 0 0 0 0 0 0 2 14 18 1 0 0 5 0 0 0 6 64 64 0 65 128 0 0 129 192 0 0 28 128 128 1 69 0 0 0 70 0 193 0 128 0 0 0 193 64 1 0 92 128 128 1 133 192 1 0 134 0 66 1 193 64 2 0 1 129 2 0 65 65 2 0 129 65 2 0 156 128 128 2 73 128 0 131 133 192 1 0 134 0 67 1 193 64 3 0 1 65 3 0 65 65 2 0 129 65 3 0 156 128 128 2 73 128 128 133 133 192 3 0 134 0 67 1 193 0 4 0 1 65 4 0 65 129 2 0 156 128 0 2 73 128 0 135 133 0 0 0 134 0 65 1 192 0 0 0 1 129 4 0 156 128 128 1 197 192 1 0 198 0 195 1 1 65 3 0 65 65 3 0 129 65 2 0 193 65 3 0 220 128 128 2 137 192 128 133 197 192 1 0 198 0 195 1 1 193 4 0 65 65 3 0 129 129 2 0 193 65 3 0 220 128 128 2 137 192 0 131 197 192 3 0 198 0 195 1 1 1 4 0 65 65 4 0 129 129 2 0 220 128 0 2 137 192 0 135 137 64 69 138 197 192 5 0 198 128 197 1 198 0 198 1 137 192 0 139 137 128 198 140 137 0 199 141 137 128 199 142 197 192 3 0 198 0 195 1 1 1 8 0 65 65 8 0 129 129 8 0 220 128 0 2 137 192 128 143 197 0 0 0 198 0 193 1 0 1 0 0 65 193 8 0 220 128 128 1 201 64 73 146 5 193 1 0 6 1 67 2 65 193 4 0 129 193 4 0 193 193 4 0 1 194 4 0 28 129 128 2 201 0 1 131 201 64 66 147 6 193 201 1 11 1 74 2 164 1 0 0 0 0 128 1 28 65 128 1 6 65 202 1 11 1 74 2 164 65 0 0 0 0 128 1 28 65 128 1 6 129 202 1 11 1 74 2 164 129 0 0 28 65 128 1 5 1 0 0 6 1 65 2 64 1 0 0 129 193 8 0 28 129 128 1 9 193 74 146 69 193 1 0 70 1 195 2 129 193 4 0 193 193 4 0 1 194 4 0 65 194 4 0 92 129 128 2 9 65 1 131 69 193 1 0 70 1 195 2 129 193 4 0 193 65 3 0 1 66 3 0 65 66 3 0 92 129 128 2 9 65 129 133 9 65 66 147 70 193 73 2 75 1 202 2 228 193 0 0 0 0 0 2 92 65 128 1 70 65 74 2 75 1 202 2 228 1 1 0 0 0 0 2 92 65 128 1 69 1 0 0 70 1 193 2 128 1 0 0 193 193 8 0 92 129 128 1 133 193 1 0 134 1 67 3 193 65 8 0 1 66 3 0 65 66 3 0 129 66 3 0 156 129 128 2 73 129 129 133 73 65 66 147 134 193 201 2 139 1 74 3 36 66 1 0 0 0 128 2 156 65 128 1 134 65 202 2 139 1 74 3 36 130 1 0 0 0 128 2 156 65 128 1 133 1 0 0 134 1 65 3 192 1 0 0 1 194 8 0 156 129 128 1 137 1 75 146 197 193 1 0 198 1 195 3 1 194 4 0 65 194 4 0 129 194 4 0 193 194 4 0 220 129 128 2 137 193 1 131 197 193 1 0 198 1 195 3 1 66 8 0 65 66 3 0 129 66 3 0 193 66 3 0 220 129 128 2 137 193 129 133 137 65 66 147 198 193 73 3 203 1 202 3 100 194 1 0 0 0 0 3 220 65 128 1 198 65 74 3 203 1 202 3 100 2 2 0 0 0 0 3 220 65 128 1 197 1 0 0 198 1 193 3 0 2 0 0 65 194 8 0 220 129 128 1 201 65 75 146 5 194 1 0 6 2 67 4 65 194 4 0 129 194 4 0 193 194 4 0 1 195 4 0 28 130 128 2 201 1 2 131 5 194 1 0 6 2 67 4 65 130 11 0 129 66 3 0 193 66 3 0 1 67 3 0 28 130 128 2 201 1 130 133 201 65 66 147 6 194 201 3 11 2 74 4 164 66 2 0 0 0 128 3 28 66 128 1 6 66 202 3 11 2 74 4 164 130 2 0 0 0 128 3 28 66 128 1 5 2 0 0 6 2 65 4 64 2 0 0 129 130 4 0 28 130 128 1 69 194 1 0 70 2 195 4 129 194 4 0 193 66 3 0 1 67 2 0 65 67 3 0 92 130 128 2 9 66 130 133 69 194 1 0 70 2 195 4 129 66 8 0 193 66 3 0 1 131 2 0 65 67 3 0 92 130 128 2 9 66 2 131 69 194 3 0 70 2 195 4 129 2 4 0 193 66 4 0 1 131 2 0 92 130 0 2 9 66 2 135 9 66 67 138 69 194 5 0 70 130 197 4 70 2 198 4 9 66 2 139 9 194 203 140 9 66 66 152 9 66 204 142 9 130 204 141 9 66 204 153 69 194 3 0 70 2 195 4 129 2 8 0 193 66 8 0 1 131 8 0 92 130 0 2 9 66 130 143 30 0 128 0 52 0 0 0 4 5 0 0 0 0 0 0 0 76 105 109 101 0 4 13 0 0 0 0 0 0 0 67 114 101 97 116 101 87 105 110 100 111 119 0 4 13 0 0 0 0 0 0 0 80 104 111 116 111 76 105 109 101 32 118 49 0 4 24 0 0 0 0 0 0 0 114 98 120 97 115 115 101 116 105 100 58 47 47 57 51 57 55 48 50 57 52 56 50 0 4 9 0 0 0 0 0 0 0 67 114 101 97 116 101 85 73 0 4 6 0 0 0 0 0 0 0 70 114 97 109 101 0 4 5 0 0 0 0 0 0 0 83 105 122 101 0 4 6 0 0 0 0 0 0 0 85 68 105 109 50 0 4 10 0 0 0 0 0 0 0 102 114 111 109 83 99 97 108 101 0 3 0 0 0 0 0 0 240 63 3 154 153 153 153 153 153 185 63 4 9 0 0 0 0 0 0 0 80 111 115 105 116 105 111 110 0 4 4 0 0 0 0 0 0 0 110 101 119 0 3 0 0 0 0 0 0 0 0 4 17 0 0 0 0 0 0 0 66 97 99 107 103 114 111 117 110 100 67 111 108 111 114 51 0 4 7 0 0 0 0 0 0 0 67 111 108 111 114 51 0 3 236 81 184 30 133 235 177 63 3 123 20 174 71 225 122 180 63 4 11 0 0 0 0 0 0 0 84 101 120 116 66 117 116 116 111 110 0 3 154 153 153 153 153 153 201 63 4 16 0 0 0 0 0 0 0 66 111 114 100 101 114 83 105 122 101 80 105 120 101 108 0 3 154 153 153 153 153 153 13 64 4 5 0 0 0 0 0 0 0 70 111 110 116 0 4 5 0 0 0 0 0 0 0 69 110 117 109 0 4 7 0 0 0 0 0 0 0 85 98 117 110 116 117 0 4 9 0 0 0 0 0 0 0 84 101 120 116 83 105 122 101 0 3 0 0 0 0 0 0 68 64 4 5 0 0 0 0 0 0 0 84 101 120 116 0 4 7 0 0 0 0 0 0 0 80 97 103 101 32 49 0 4 11 0 0 0 0 0 0 0 84 101 120 116 83 99 97 108 101 100 0 1 1 4 11 0 0 0 0 0 0 0 84 101 120 116 67 111 108 111 114 51 0 3 51 51 51 51 51 51 211 63 3 154 153 153 153 153 153 217 63 3 0 0 0 0 0 0 224 63 4 12 0 0 0 0 0 0 0 73 109 97 103 101 66 117 116 116 111 110 0 4 6 0 0 0 0 0 0 0 73 109 97 103 101 0 4 43 0 0 0 0 0 0 0 104 116 116 112 58 47 47 119 119 119 46 114 111 98 108 111 120 46 99 111 109 47 97 115 115 101 116 47 63 105 100 61 56 52 50 53 48 54 57 55 49 56 0 4 7 0 0 0 0 0 0 0 90 73 110 100 101 120 0 4 11 0 0 0 0 0 0 0 77 111 117 115 101 69 110 116 101 114 0 4 8 0 0 0 0 0 0 0 67 111 110 110 101 99 116 0 4 11 0 0 0 0 0 0 0 77 111 117 115 101 76 101 97 118 101 0 4 18 0 0 0 0 0 0 0 77 111 117 115 101 66 117 116 116 111 110 49 67 108 105 99 107 0 4 43 0 0 0 0 0 0 0 104 116 116 112 58 47 47 119 119 119 46 114 111 98 108 111 120 46 99 111 109 47 97 115 115 101 116 47 63 105 100 61 56 51 52 53 56 53 56 49 49 52 0 4 43 0 0 0 0 0 0 0 104 116 116 112 58 47 47 119 119 119 46 114 111 98 108 111 120 46 99 111 109 47 97 115 115 101 116 47 63 105 100 61 56 52 53 48 54 48 49 51 53 49 0 4 43 0 0 0 0 0 0 0 104 116 116 112 58 47 47 119 119 119 46 114 111 98 108 111 120 46 99 111 109 47 97 115 115 101 116 47 63 105 100 61 54 48 55 53 51 57 53 56 52 54 0 3 51 51 51 51 51 51 227 63 3 0 0 0 0 0 0 54 64 4 23 0 0 0 0 0 0 0 66 97 99 107 103 114 111 117 110 100 84 114 97 110 115 112 97 114 101 110 99 121 0 1 0 4 11 0 0 0 0 0 0 0 77 111 114 101 32 83 111 111 110 33 0 4 7 0 0 0 0 0 0 0 65 99 116 105 118 101 0 11 0 0 0 0 0 0 0 0 0 0 0 26 0 0 0 29 0 0 0 1 0 0 6 12 0 0 0 4 0 0 0 69 64 0 0 70 128 192 0 129 192 0 0 193 192 0 0 1 193 0 0 65 193 0 0 92 128 128 2 9 64 0 128 4 0 0 0 9 64 65 130 30 0 128 0 6 0 0 0 4 5 0 0 0 0 0 0 0 83 105 122 101 0 4 6 0 0 0 0 0 0 0 85 68 105 109 50 0 4 4 0 0 0 0 0 0 0 110 101 119 0 3 31 133 235 81 184 30 213 63 4 7 0 0 0 0 0 0 0 90 73 110 100 101 120 0 3 0 0 0 0 0 0 0 64 0 0 0 0 12 0 0 0 27 0 0 0 27 0 0 0 27 0 0 0 27 0 0 0 27 0 0 0 27 0 0 0 27 0 0 0 27 0 0 0 27 0 0 0 28 0 0 0 28 0 0 0 29 0 0 0 0 0 0 0 1 0 0 0 7 0 0 0 0 0 0 0 73 109 97 103 101 49 0 0 0 0 0 0 0 0 0 31 0 0 0 34 0 0 0 1 0 0 6 12 0 0 0 4 0 0 0 69 64 0 0 70 128 192 0 129 192 0 0 193 192 0 0 1 193 0 0 65 193 0 0 92 128 128 2 9 64 0 128 4 0 0 0 9 64 65 130 30 0 128 0 6 0 0 0 4 5 0 0 0 0 0 0 0 83 105 122 101 0 4 6 0 0 0 0 0 0 0 85 68 105 109 50 0 4 4 0 0 0 0 0 0 0 110 101 119 0 3 154 153 153 153 153 153 201 63 4 7 0 0 0 0 0 0 0 90 73 110 100 101 120 0 3 0 0 0 0 0 0 240 63 0 0 0 0 12 0 0 0 32 0 0 0 32 0 0 0 32 0 0 0 32 0 0 0 32 0 0 0 32 0 0 0 32 0 0 0 32 0 0 0 32 0 0 0 33 0 0 0 33 0 0 0 34 0 0 0 0 0 0 0 1 0 0 0 7 0 0 0 0 0 0 0 73 109 97 103 101 49 0 0 0 0 0 0 0 0 0 36 0 0 0 38 0 0 0 0 0 0 2 1 0 0 0 30 0 128 0 0 0 0 0 0 0 0 0 1 0 0 0 38 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 46 0 0 0 49 0 0 0 1 0 0 6 12 0 0 0 4 0 0 0 69 64 0 0 70 128 192 0 129 192 0 0 193 192 0 0 1 193 0 0 65 193 0 0 92 128 128 2 9 64 0 128 4 0 0 0 9 64 65 130 30 0 128 0 6 0 0 0 4 5 0 0 0 0 0 0 0 83 105 122 101 0 4 6 0 0 0 0 0 0 0 85 68 105 109 50 0 4 4 0 0 0 0 0 0 0 110 101 119 0 3 31 133 235 81 184 30 213 63 4 7 0 0 0 0 0 0 0 90 73 110 100 101 120 0 3 0 0 0 0 0 0 0 64 0 0 0 0 12 0 0 0 47 0 0 0 47 0 0 0 47 0 0 0 47 0 0 0 47 0 0 0 47 0 0 0 47 0 0 0 47 0 0 0 47 0 0 0 48 0 0 0 48 0 0 0 49 0 0 0 0 0 0 0 1 0 0 0 7 0 0 0 0 0 0 0 73 109 97 103 101 50 0 0 0 0 0 0 0 0 0 51 0 0 0 54 0 0 0 1 0 0 6 12 0 0 0 4 0 0 0 69 64 0 0 70 128 192 0 129 192 0 0 193 192 0 0 1 193 0 0 65 193 0 0 92 128 128 2 9 64 0 128 4 0 0 0 9 64 65 130 30 0 128 0 6 0 0 0 4 5 0 0 0 0 0 0 0 83 105 122 101 0 4 6 0 0 0 0 0 0 0 85 68 105 109 50 0 4 4 0 0 0 0 0 0 0 110 101 119 0 3 154 153 153 153 153 153 201 63 4 7 0 0 0 0 0 0 0 90 73 110 100 101 120 0 3 0 0 0 0 0 0 240 63 0 0 0 0 12 0 0 0 52 0 0 0 52 0 0 0 52 0 0 0 52 0 0 0 52 0 0 0 52 0 0 0 52 0 0 0 52 0 0 0 52 0 0 0 53 0 0 0 53 0 0 0 54 0 0 0 0 0 0 0 1 0 0 0 7 0 0 0 0 0 0 0 73 109 97 103 101 50 0 0 0 0 0 0 0 0 0 61 0 0 0 64 0 0 0 1 0 0 6 12 0 0 0 4 0 0 0 69 64 0 0 70 128 192 0 129 192 0 0 193 192 0 0 1 193 0 0 65 193 0 0 92 128 128 2 9 64 0 128 4 0 0 0 9 64 65 130 30 0 128 0 6 0 0 0 4 5 0 0 0 0 0 0 0 83 105 122 101 0 4 6 0 0 0 0 0 0 0 85 68 105 109 50 0 4 4 0 0 0 0 0 0 0 110 101 119 0 3 31 133 235 81 184 30 213 63 4 7 0 0 0 0 0 0 0 90 73 110 100 101 120 0 3 0 0 0 0 0 0 0 64 0 0 0 0 12 0 0 0 62 0 0 0 62 0 0 0 62 0 0 0 62 0 0 0 62 0 0 0 62 0 0 0 62 0 0 0 62 0 0 0 62 0 0 0 63 0 0 0 63 0 0 0 64 0 0 0 0 0 0 0 1 0 0 0 7 0 0 0 0 0 0 0 73 109 97 103 101 51 0 0 0 0 0 0 0 0 0 66 0 0 0 69 0 0 0 1 0 0 6 12 0 0 0 4 0 0 0 69 64 0 0 70 128 192 0 129 192 0 0 193 192 0 0 1 193 0 0 65 193 0 0 92 128 128 2 9 64 0 128 4 0 0 0 9 64 65 130 30 0 128 0 6 0 0 0 4 5 0 0 0 0 0 0 0 83 105 122 101 0 4 6 0 0 0 0 0 0 0 85 68 105 109 50 0 4 4 0 0 0 0 0 0 0 110 101 119 0 3 154 153 153 153 153 153 201 63 4 7 0 0 0 0 0 0 0 90 73 110 100 101 120 0 3 0 0 0 0 0 0 240 63 0 0 0 0 12 0 0 0 67 0 0 0 67 0 0 0 67 0 0 0 67 0 0 0 67 0 0 0 67 0 0 0 67 0 0 0 67 0 0 0 67 0 0 0 68 0 0 0 68 0 0 0 69 0 0 0 0 0 0 0 1 0 0 0 7 0 0 0 0 0 0 0 73 109 97 103 101 51 0 0 0 0 0 0 0 0 0 78 0 0 0 81 0 0 0 1 0 0 6 12 0 0 0 4 0 0 0 69 64 0 0 70 128 192 0 129 192 0 0 193 192 0 0 1 193 0 0 65 193 0 0 92 128 128 2 9 64 0 128 4 0 0 0 9 64 65 130 30 0 128 0 6 0 0 0 4 5 0 0 0 0 0 0 0 83 105 122 101 0 4 6 0 0 0 0 0 0 0 85 68 105 109 50 0 4 4 0 0 0 0 0 0 0 110 101 119 0 3 31 133 235 81 184 30 213 63 4 7 0 0 0 0 0 0 0 90 73 110 100 101 120 0 3 0 0 0 0 0 0 0 64 0 0 0 0 12 0 0 0 79 0 0 0 79 0 0 0 79 0 0 0 79 0 0 0 79 0 0 0 79 0 0 0 79 0 0 0 79 0 0 0 79 0 0 0 80 0 0 0 80 0 0 0 81 0 0 0 0 0 0 0 1 0 0 0 7 0 0 0 0 0 0 0 73 109 97 103 101 52 0 0 0 0 0 0 0 0 0 83 0 0 0 86 0 0 0 1 0 0 6 12 0 0 0 4 0 0 0 69 64 0 0 70 128 192 0 129 192 0 0 193 192 0 0 1 193 0 0 65 193 0 0 92 128 128 2 9 64 0 128 4 0 0 0 9 64 65 130 30 0 128 0 6 0 0 0 4 5 0 0 0 0 0 0 0 83 105 122 101 0 4 6 0 0 0 0 0 0 0 85 68 105 109 50 0 4 4 0 0 0 0 0 0 0 110 101 119 0 3 154 153 153 153 153 153 201 63 4 7 0 0 0 0 0 0 0 90 73 110 100 101 120 0 3 0 0 0 0 0 0 240 63 0 0 0 0 12 0 0 0 84 0 0 0 84 0 0 0 84 0 0 0 84 0 0 0 84 0 0 0 84 0 0 0 84 0 0 0 84 0 0 0 84 0 0 0 85 0 0 0 85 0 0 0 86 0 0 0 0 0 0 0 1 0 0 0 7 0 0 0 0 0 0 0 73 109 97 103 101 52 0 0 0 0 0 0 0 0 0 95 0 0 0 98 0 0 0 1 0 0 6 12 0 0 0 4 0 0 0 69 64 0 0 70 128 192 0 129 192 0 0 193 192 0 0 1 193 0 0 65 193 0 0 92 128 128 2 9 64 0 128 4 0 0 0 9 64 65 130 30 0 128 0 6 0 0 0 4 5 0 0 0 0 0 0 0 83 105 122 101 0 4 6 0 0 0 0 0 0 0 85 68 105 109 50 0 4 4 0 0 0 0 0 0 0 110 101 119 0 3 31 133 235 81 184 30 213 63 4 7 0 0 0 0 0 0 0 90 73 110 100 101 120 0 3 0 0 0 0 0 0 0 64 0 0 0 0 12 0 0 0 96 0 0 0 96 0 0 0 96 0 0 0 96 0 0 0 96 0 0 0 96 0 0 0 96 0 0 0 96 0 0 0 96 0 0 0 97 0 0 0 97 0 0 0 98 0 0 0 0 0 0 0 1 0 0 0 7 0 0 0 0 0 0 0 73 109 97 103 101 53 0 0 0 0 0 0 0 0 0 100 0 0 0 103 0 0 0 1 0 0 6 12 0 0 0 4 0 0 0 69 64 0 0 70 128 192 0 129 192 0 0 193 192 0 0 1 193 0 0 65 193 0 0 92 128 128 2 9 64 0 128 4 0 0 0 9 64 65 130 30 0 128 0 6 0 0 0 4 5 0 0 0 0 0 0 0 83 105 122 101 0 4 6 0 0 0 0 0 0 0 85 68 105 109 50 0 4 4 0 0 0 0 0 0 0 110 101 119 0 3 154 153 153 153 153 153 201 63 4 7 0 0 0 0 0 0 0 90 73 110 100 101 120 0 3 0 0 0 0 0 0 240 63 0 0 0 0 12 0 0 0 101 0 0 0 101 0 0 0 101 0 0 0 101 0 0 0 101 0 0 0 101 0 0 0 101 0 0 0 101 0 0 0 101 0 0 0 102 0 0 0 102 0 0 0 103 0 0 0 0 0 0 0 1 0 0 0 7 0 0 0 0 0 0 0 73 109 97 103 101 53 0 18 1 0 0 3 0 0 0 3 0 0 0 3 0 0 0 3 0 0 0 3 0 0 0 5 0 0 0 5 0 0 0 5 0 0 0 5 0 0 0 5 0 0 0 6 0 0 0 6 0 0 0 6 0 0 0 6 0 0 0 6 0 0 0 6 0 0 0 6 0 0 0 6 0 0 0 7 0 0 0 7 0 0 0 7 0 0 0 7 0 0 0 7 0 0 0 7 0 0 0 7 0 0 0 7 0 0 0 8 0 0 0 8 0 0 0 8 0 0 0 8 0 0 0 8 0 0 0 8 0 0 0 8 0 0 0 10 0 0 0 10 0 0 0 10 0 0 0 10 0 0 0 10 0 0 0 11 0 0 0 11 0 0 0 11 0 0 0 11 0 0 0 11 0 0 0 11 0 0 0 11 0 0 0 11 0 0 0 12 0 0 0 12 0 0 0 12 0 0 0 12 0 0 0 12 0 0 0 12 0 0 0 12 0 0 0 12 0 0 0 13 0 0 0 13 0 0 0 13 0 0 0 13 0 0 0 13 0 0 0 13 0 0 0 13 0 0 0 14 0 0 0 15 0 0 0 15 0 0 0 15 0 0 0 15 0 0 0 16 0 0 0 17 0 0 0 18 0 0 0 19 0 0 0 19 0 0 0 19 0 0 0 19 0 0 0 19 0 0 0 19 0 0 0 19 0 0 0 21 0 0 0 21 0 0 0 21 0 0 0 21 0 0 0 21 0 0 0 22 0 0 0 23 0 0 0 23 0 0 0 23 0 0 0 23 0 0 0 23 0 0 0 23 0 0 0 23 0 0 0 23 0 0 0 24 0 0 0 26 0 0 0 26 0 0 0 29 0 0 0 29 0 0 0 26 0 0 0 31 0 0 0 31 0 0 0 34 0 0 0 34 0 0 0 31 0 0 0 36 0 0 0 36 0 0 0 38 0 0 0 36 0 0 0 40 0 0 0 40 0 0 0 40 0 0 0 40 0 0 0 40 0 0 0 41 0 0 0 42 0 0 0 42 0 0 0 42 0 0 0 42 0 0 0 42 0 0 0 42 0 0 0 42 0 0 0 42 0 0 0 43 0 0 0 43 0 0 0 43 0 0 0 43 0 0 0 43 0 0 0 43 0 0 0 43 0 0 0 43 0 0 0 44 0 0 0 46 0 0 0 46 0 0 0 49 0 0 0 49 0 0 0 46 0 0 0 51 0 0 0 51 0 0 0 54 0 0 0 54 0 0 0 51 0 0 0 56 0 0 0 56 0 0 0 56 0 0 0 56 0 0 0 56 0 0 0 58 0 0 0 58 0 0 0 58 0 0 0 58 0 0 0 58 0 0 0 58 0 0 0 58 0 0 0 58 0 0 0 59 0 0 0 61 0 0 0 61 0 0 0 64 0 0 0 64 0 0 0 61 0 0 0 66 0 0 0 66 0 0 0 69 0 0 0 69 0 0 0 66 0 0 0 72 0 0 0 72 0 0 0 72 0 0 0 72 0 0 0 72 0 0 0 73 0 0 0 74 0 0 0 74 0 0 0 74 0 0 0 74 0 0 0 74 0 0 0 74 0 0 0 74 0 0 0 74 0 0 0 75 0 0 0 75 0 0 0 75 0 0 0 75 0 0 0 75 0 0 0 75 0 0 0 75 0 0 0 75 0 0 0 76 0 0 0 78 0 0 0 78 0 0 0 81 0 0 0 81 0 0 0 78 0 0 0 83 0 0 0 83 0 0 0 86 0 0 0 86 0 0 0 83 0 0 0 89 0 0 0 89 0 0 0 89 0 0 0 89 0 0 0 89 0 0 0 90 0 0 0 91 0 0 0 91 0 0 0 91 0 0 0 91 0 0 0 91 0 0 0 91 0 0 0 91 0 0 0 91 0 0 0 92 0 0 0 92 0 0 0 92 0 0 0 92 0 0 0 92 0 0 0 92 0 0 0 92 0 0 0 92 0 0 0 93 0 0 0 95 0 0 0 95 0 0 0 98 0 0 0 98 0 0 0 95 0 0 0 100 0 0 0 100 0 0 0 103 0 0 0 103 0 0 0 100 0 0 0 105 0 0 0 105 0 0 0 105 0 0 0 105 0 0 0 105 0 0 0 106 0 0 0 106 0 0 0 106 0 0 0 106 0 0 0 106 0 0 0 106 0 0 0 106 0 0 0 106 0 0 0 107 0 0 0 107 0 0 0 107 0 0 0 107 0 0 0 107 0 0 0 107 0 0 0 107 0 0 0 107 0 0 0 108 0 0 0 108 0 0 0 108 0 0 0 108 0 0 0 108 0 0 0 108 0 0 0 108 0 0 0 109 0 0 0 110 0 0 0 110 0 0 0 110 0 0 0 110 0 0 0 111 0 0 0 112 0 0 0 113 0 0 0 114 0 0 0 115 0 0 0 117 0 0 0 117 0 0 0 117 0 0 0 117 0 0 0 117 0 0 0 117 0 0 0 117 0 0 0 117 0 0 0 9 0 0 0 4 0 0 0 0 0 0 0 97 112 112 0 5 0 0 0 17 1 0 0 4 0 0 0 0 0 0 0 98 97 114 0 10 0 0 0 17 1 0 0 11 0 0 0 0 0 0 0 72 111 109 101 66 117 116 116 111 110 0 38 0 0 0 17 1 0 0 7 0 0 0 0 0 0 0 73 109 97 103 101 49 0 81 0 0 0 17 1 0 0 7 0 0 0 0 0 0 0 73 109 97 103 101 50 0 110 0 0 0 17 1 0 0 7 0 0 0 0 0 0 0 73 109 97 103 101 51 0 143 0 0 0 17 1 0 0 7 0 0 0 0 0 0 0 73 109 97 103 101 52 0 167 0 0 0 17 1 0 0 7 0 0 0 0 0 0 0 73 109 97 103 101 53 0 200 0 0 0 17 1 0 0 12 0 0 0 0 0 0 0 72 111 109 101 66 117 116 116 111 110 50 0 233 0 0 0 17 1 0 0 0 0 0 0 