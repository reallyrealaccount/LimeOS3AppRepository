76 69 70 0 0 0 0 0 1 0 0 0 0 0 0 0 57 66 105 116 66 121 116 101 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 101 54 49 51 50 54 48 49 102 55 99 52 101 99 50 56 56 100 48 99 97 56 55 55 56 100 102 97 102 54 51 50 53 102 56 51 55 53 101 52 57 53 54 49 48 53 51 56 54 57 50 55 100 97 51 101 55 54 99 48 56 55 52 48 27 76 117 97 81 0 1 4 8 4 8 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 2 20 94 0 0 0 5 64 0 0 65 128 0 0 28 128 0 1 7 0 0 0 5 64 0 0 65 0 1 0 28 128 0 1 7 192 0 0 5 64 0 0 65 128 1 0 28 128 0 1 7 64 1 0 5 64 0 0 65 0 2 0 28 128 0 1 7 192 1 0 5 64 0 0 65 128 2 0 130 0 128 0 28 128 128 1 7 64 2 0 10 0 1 0 9 64 67 134 9 192 67 135 9 64 68 136 9 192 68 137 7 192 2 0 10 0 0 9 65 64 5 0 129 128 5 0 193 192 5 0 1 1 6 0 65 65 6 0 129 129 6 0 193 193 6 0 1 2 7 0 65 66 7 0 129 130 7 0 193 194 7 0 1 3 8 0 65 67 8 0 129 131 8 0 193 195 8 0 1 4 9 0 65 68 9 0 129 132 9 0 193 196 9 0 34 64 128 9 7 0 5 0 1 64 10 0 7 0 10 0 1 192 10 0 7 128 10 0 1 64 11 0 7 0 11 0 1 192 11 0 7 128 11 0 5 0 0 0 6 0 76 0 65 64 12 0 28 64 0 1 5 192 12 0 69 128 10 0 129 0 13 0 197 0 11 0 28 128 0 2 7 128 12 0 2 0 128 0 66 0 0 0 164 0 0 0 135 64 13 0 164 64 0 0 135 0 3 0 164 128 0 0 135 128 3 0 164 192 0 0 135 128 13 0 164 0 1 0 135 192 13 0 164 64 1 0 135 0 14 0 164 128 1 0 135 64 14 0 164 192 1 0 0 0 128 0 135 128 14 0 164 0 2 0 135 192 14 0 164 64 2 0 0 0 0 0 135 0 15 0 133 0 15 0 156 64 128 0 30 0 128 0 61 0 0 0 4 5 0 0 0 0 0 0 0 107 114 110 108 0 4 8 0 0 0 0 0 0 0 108 111 97 100 108 105 98 0 4 11 0 0 0 0 0 0 0 76 105 109 101 75 101 114 110 101 108 0 4 3 0 0 0 0 0 0 0 97 102 0 4 17 0 0 0 0 0 0 0 76 105 109 101 65 112 112 70 114 97 109 101 119 111 114 107 0 4 4 0 0 0 0 0 0 0 101 120 112 0 4 13 0 0 0 0 0 0 0 76 105 109 101 69 120 112 108 111 114 101 114 0 4 5 0 0 0 0 0 0 0 110 111 116 105 0 4 18 0 0 0 0 0 0 0 76 105 109 101 78 111 116 105 102 105 99 97 116 105 111 110 115 0 4 11 0 0 0 0 0 0 0 108 111 97 100 115 116 114 105 110 103 0 4 11 0 0 0 0 0 0 0 76 111 97 100 115 116 114 105 110 103 0 4 7 0 0 0 0 0 0 0 101 114 114 111 114 115 0 4 8 0 0 0 0 0 0 0 69 82 82 95 53 48 51 0 4 127 0 0 0 0 0 0 0 60 98 62 69 82 82 95 53 48 51 60 47 98 62 32 124 32 80 114 111 119 115 101 114 32 105 115 32 99 117 114 114 101 110 116 108 121 32 110 111 116 32 97 118 97 105 108 97 98 108 101 33 32 84 104 105 115 32 105 115 32 101 105 116 104 101 114 32 100 117 101 32 116 111 32 109 97 105 110 116 101 110 97 110 99 101 32 111 114 32 97 32 115 104 117 116 100 111 119 110 46 32 80 108 101 97 115 101 32 99 104 101 99 107 32 98 97 99 107 32 108 97 116 101 114 46 0 4 12 0 0 0 0 0 0 0 69 82 82 95 87 69 66 95 52 48 52 0 4 114 0 0 0 0 0 0 0 60 98 62 69 82 82 95 87 69 66 95 52 48 52 60 47 98 62 32 124 32 84 104 101 32 114 101 113 117 101 115 116 101 100 32 115 105 116 101 32 119 97 115 32 110 111 116 32 102 111 117 110 100 46 32 80 108 101 97 115 101 32 99 104 101 99 107 32 121 111 117 114 32 115 112 101 108 108 105 110 103 44 32 97 110 100 32 109 97 107 101 32 115 117 114 101 32 116 104 101 32 115 105 116 101 32 101 120 105 115 116 115 33 0 4 12 0 0 0 0 0 0 0 69 82 82 95 87 69 66 95 52 48 48 0 4 100 0 0 0 0 0 0 0 60 98 62 69 82 82 95 87 69 66 95 52 48 48 60 47 98 62 32 124 32 84 104 101 32 98 114 111 119 115 101 114 32 119 97 115 32 117 110 97 98 108 101 32 116 111 32 114 101 99 105 101 118 101 32 100 97 116 97 46 32 84 104 105 115 32 109 97 121 32 98 101 32 97 32 110 101 116 119 111 114 107 32 111 114 32 82 111 98 108 111 120 32 105 115 115 117 101 46 0 4 12 0 0 0 0 0 0 0 69 82 82 95 87 69 66 95 52 48 49 0 4 93 0 0 0 0 0 0 0 60 98 62 69 82 82 95 87 69 66 95 52 48 49 60 47 98 62 32 124 32 89 111 117 114 32 99 108 105 101 110 116 32 100 111 101 115 32 110 111 116 32 104 97 118 101 32 116 104 101 32 112 114 111 112 101 114 32 112 101 114 109 105 115 115 105 111 110 115 32 116 111 32 118 105 101 119 32 116 104 105 115 32 114 101 115 111 117 114 99 101 46 0 4 10 0 0 0 0 0 0 0 102 105 108 101 110 97 109 101 115 0 4 4 0 0 0 0 0 0 0 76 105 98 0 4 11 0 0 0 0 0 0 0 77 111 100 117 108 101 77 97 105 110 0 4 11 0 0 0 0 0 0 0 71 105 116 76 105 98 114 97 114 121 0 4 12 0 0 0 0 0 0 0 80 114 111 119 115 101 114 77 97 105 110 0 4 10 0 0 0 0 0 0 0 80 114 111 119 115 101 114 83 72 0 4 8 0 0 0 0 0 0 0 69 78 67 108 111 97 100 0 4 8 0 0 0 0 0 0 0 69 84 72 108 111 97 100 0 4 6 0 0 0 0 0 0 0 83 72 115 101 116 0 4 9 0 0 0 0 0 0 0 72 71 121 103 55 54 71 84 0 4 7 0 0 0 0 0 0 0 83 101 116 80 111 115 0 4 7 0 0 0 0 0 0 0 71 101 116 80 111 115 0 4 6 0 0 0 0 0 0 0 87 101 98 71 76 0 4 8 0 0 0 0 0 0 0 76 105 109 101 78 69 84 0 4 13 0 0 0 0 0 0 0 80 114 111 119 115 101 114 85 115 101 114 115 0 4 23 0 0 0 0 0 0 0 108 111 99 97 108 58 47 47 49 50 55 46 48 46 48 46 49 58 53 53 48 48 0 4 7 0 0 0 0 0 0 0 47 73 110 105 116 47 0 4 4 0 0 0 0 0 0 0 82 101 103 0 4 13 0 0 0 0 0 0 0 83 105 116 101 82 101 103 105 115 116 114 121 0 4 8 0 0 0 0 0 0 0 87 101 98 70 117 110 99 0 4 15 0 0 0 0 0 0 0 115 105 116 101 115 85 82 76 112 114 101 102 105 120 0 4 68 0 0 0 0 0 0 0 104 116 116 112 115 58 47 47 114 97 119 46 103 105 116 104 117 98 117 115 101 114 99 111 110 116 101 110 116 46 99 111 109 47 66 97 114 114 97 99 117 100 97 76 97 107 101 47 76 105 109 101 78 101 116 47 109 97 105 110 47 115 105 116 101 115 47 0 4 5 0 0 0 0 0 0 0 110 97 109 101 0 4 38 0 0 0 0 0 0 0 80 82 79 87 83 69 82 32 45 32 73 110 116 101 114 110 101 116 32 66 114 111 119 115 101 114 32 102 111 114 32 76 105 109 101 79 83 0 4 7 0 0 0 0 0 0 0 108 111 103 111 73 100 0 4 25 0 0 0 0 0 0 0 114 98 120 97 115 115 101 116 105 100 58 47 47 49 49 51 54 54 50 51 53 53 51 51 0 4 10 0 0 0 0 0 0 0 108 111 103 111 73 100 82 97 119 0 3 0 0 104 236 215 43 5 66 4 12 0 0 0 0 0 0 0 65 108 108 111 99 97 116 101 82 97 109 0 3 0 0 0 0 0 128 65 64 4 4 0 0 0 0 0 0 0 97 112 112 0 4 10 0 0 0 0 0 0 0 99 114 101 97 116 101 97 112 112 0 3 0 0 0 0 0 0 240 63 4 12 0 0 0 0 0 0 0 101 114 114 111 114 95 102 114 97 109 101 0 4 10 0 0 0 0 0 0 0 83 101 108 101 99 116 84 97 98 0 4 7 0 0 0 0 0 0 0 78 101 119 84 97 98 0 4 21 0 0 0 0 0 0 0 76 111 111 112 84 101 120 116 84 114 97 110 115 112 97 114 101 110 99 121 0 4 11 0 0 0 0 0 0 0 67 104 97 110 103 101 84 101 120 116 0 4 7 0 0 0 0 0 0 0 83 101 97 114 99 104 0 4 5 0 0 0 0 0 0 0 73 110 105 116 0 4 5 0 0 0 0 0 0 0 108 111 97 100 0 10 0 0 0 0 0 0 0 0 0 0 0 29 0 0 0 51 0 0 0 0 0 0 4 89 0 0 0 5 64 0 0 65 128 0 0 133 192 0 0 28 128 128 1 7 0 0 0 5 0 0 0 69 64 1 0 70 128 193 0 129 192 1 0 193 192 1 0 92 128 128 1 9 64 0 130 5 64 0 0 65 64 2 0 133 0 0 0 28 128 128 1 7 0 2 0 5 0 2 0 69 64 1 0 70 128 193 0 129 128 2 0 193 192 2 0 92 128 128 1 9 64 0 130 5 0 2 0 69 64 1 0 70 128 193 0 129 64 3 0 193 128 3 0 92 128 128 1 9 64 0 134 5 0 2 0 9 0 196 135 5 0 2 0 69 128 4 0 70 64 196 0 70 192 196 0 9 64 128 136 5 0 2 0 69 128 4 0 70 0 197 0 70 64 197 0 9 64 0 138 5 0 2 0 9 192 69 139 5 0 2 0 9 192 65 140 5 64 0 0 65 64 2 0 133 0 0 0 28 128 128 1 7 64 6 0 5 64 6 0 9 192 70 141 5 64 6 0 69 64 1 0 70 128 193 0 129 64 3 0 193 0 7 0 92 128 128 1 9 64 0 134 5 64 6 0 69 64 1 0 70 128 193 0 129 64 7 0 193 128 7 0 92 128 128 1 9 64 0 130 5 64 6 0 69 128 4 0 70 64 196 0 70 192 196 0 9 64 128 136 5 64 6 0 9 192 197 143 5 64 6 0 9 0 200 135 5 64 6 0 69 128 4 0 70 0 197 0 70 64 197 0 9 64 0 138 5 64 6 0 9 192 69 139 5 64 6 0 9 192 65 140 5 0 0 0 30 0 0 1 30 0 128 0 33 0 0 0 4 6 0 0 0 0 0 0 0 102 114 97 109 101 0 4 4 0 0 0 0 0 0 0 110 101 119 0 4 6 0 0 0 0 0 0 0 70 114 97 109 101 0 4 4 0 0 0 0 0 0 0 97 112 112 0 4 5 0 0 0 0 0 0 0 83 105 122 101 0 4 6 0 0 0 0 0 0 0 85 68 105 109 50 0 4 10 0 0 0 0 0 0 0 102 114 111 109 83 99 97 108 101 0 3 0 0 0 0 0 0 240 63 4 5 0 0 0 0 0 0 0 116 101 120 116 0 4 10 0 0 0 0 0 0 0 84 101 120 116 76 97 98 101 108 0 3 0 0 0 0 0 0 232 63 3 51 51 51 51 51 51 195 63 4 9 0 0 0 0 0 0 0 80 111 115 105 116 105 111 110 0 3 154 153 153 153 153 153 185 63 3 0 0 0 0 0 0 208 63 4 5 0 0 0 0 0 0 0 84 101 120 116 0 4 3 0 0 0 0 0 0 0 58 40 0 4 5 0 0 0 0 0 0 0 70 111 110 116 0 4 5 0 0 0 0 0 0 0 69 110 117 109 0 4 5 0 0 0 0 0 0 0 67 111 100 101 0 4 15 0 0 0 0 0 0 0 84 101 120 116 88 65 108 105 103 110 109 101 110 116 0 4 5 0 0 0 0 0 0 0 76 101 102 116 0 4 11 0 0 0 0 0 0 0 84 101 120 116 83 99 97 108 101 100 0 1 1 4 23 0 0 0 0 0 0 0 66 97 99 107 103 114 111 117 110 100 84 114 97 110 115 112 97 114 101 110 99 121 0 4 10 0 0 0 0 0 0 0 101 114 114 111 114 99 111 100 101 0 4 5 0 0 0 0 0 0 0 78 97 109 101 0 4 10 0 0 0 0 0 0 0 69 114 114 111 114 84 101 120 116 0 3 205 204 204 204 204 204 220 63 3 51 51 51 51 51 51 235 63 3 154 153 153 153 153 153 201 63 4 9 0 0 0 0 0 0 0 82 105 99 104 84 101 120 116 0 4 27 0 0 0 0 0 0 0 65 110 32 117 110 107 110 111 119 110 32 101 114 114 111 114 32 111 99 99 117 114 114 101 100 46 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 53 0 0 0 57 0 0 0 0 1 0 3 11 0 0 0 75 0 64 0 92 64 0 1 69 128 0 0 92 128 128 0 71 64 0 0 69 64 0 0 70 192 192 0 133 64 1 0 134 128 65 1 73 128 0 130 30 0 128 0 7 0 0 0 4 8 0 0 0 0 0 0 0 68 101 115 116 114 111 121 0 4 5 0 0 0 0 0 0 0 101 114 114 102 0 4 12 0 0 0 0 0 0 0 101 114 114 111 114 95 102 114 97 109 101 0 4 10 0 0 0 0 0 0 0 69 114 114 111 114 84 101 120 116 0 4 5 0 0 0 0 0 0 0 84 101 120 116 0 4 7 0 0 0 0 0 0 0 101 114 114 111 114 115 0 4 8 0 0 0 0 0 0 0 69 82 82 95 53 48 51 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 59 0 0 0 65 0 0 0 0 1 0 3 15 0 0 0 70 64 64 0 71 0 0 0 70 192 64 0 71 128 0 0 75 0 65 0 92 64 0 1 69 128 1 0 92 128 128 0 71 64 1 0 69 64 1 0 70 192 193 0 133 64 2 0 134 128 66 1 73 128 0 132 30 0 128 0 11 0 0 0 4 4 0 0 0 0 0 0 0 112 111 115 0 4 9 0 0 0 0 0 0 0 80 111 115 105 116 105 111 110 0 4 5 0 0 0 0 0 0 0 115 105 122 101 0 4 5 0 0 0 0 0 0 0 83 105 122 101 0 4 8 0 0 0 0 0 0 0 68 101 115 116 114 111 121 0 4 5 0 0 0 0 0 0 0 101 114 114 102 0 4 12 0 0 0 0 0 0 0 101 114 114 111 114 95 102 114 97 109 101 0 4 10 0 0 0 0 0 0 0 69 114 114 111 114 84 101 120 116 0 4 5 0 0 0 0 0 0 0 84 101 120 116 0 4 7 0 0 0 0 0 0 0 101 114 114 111 114 115 0 4 12 0 0 0 0 0 0 0 69 82 82 95 87 69 66 95 52 48 52 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 67 0 0 0 69 0 0 0 0 1 0 2 1 0 0 0 30 0 128 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 71 0 0 0 89 0 0 0 0 1 0 7 52 0 0 0 69 0 0 0 129 64 0 0 92 128 0 1 133 0 0 0 193 128 0 0 0 1 128 0 156 128 128 1 197 0 1 0 198 64 193 1 1 129 1 0 65 193 1 0 129 1 2 0 220 128 0 2 73 192 128 129 197 128 2 0 198 192 194 1 1 1 3 0 65 65 3 0 220 128 128 1 73 192 128 132 203 128 195 0 65 193 3 0 130 1 0 0 220 64 0 2 197 0 1 0 198 64 193 1 1 65 4 0 65 65 4 0 129 65 4 0 220 128 0 2 137 192 0 136 73 192 68 137 137 0 69 137 197 128 2 0 198 192 194 1 1 129 5 0 65 193 5 0 220 128 128 1 137 192 128 138 197 128 2 0 198 192 194 1 1 1 6 0 65 65 3 0 220 128 128 1 137 192 128 132 137 64 195 140 137 192 70 141 137 64 71 142 137 192 71 143 73 192 69 144 94 0 0 1 30 0 128 0 33 0 0 0 4 4 0 0 0 0 0 0 0 110 101 119 0 4 11 0 0 0 0 0 0 0 84 101 120 116 66 117 116 116 111 110 0 4 10 0 0 0 0 0 0 0 84 101 120 116 76 97 98 101 108 0 4 17 0 0 0 0 0 0 0 66 97 99 107 103 114 111 117 110 100 67 111 108 111 114 51 0 4 7 0 0 0 0 0 0 0 67 111 108 111 114 51 0 4 8 0 0 0 0 0 0 0 102 114 111 109 82 71 66 0 3 0 0 0 0 0 0 59 64 3 0 0 0 0 0 0 73 64 3 0 0 0 0 0 0 95 64 4 5 0 0 0 0 0 0 0 83 105 122 101 0 4 6 0 0 0 0 0 0 0 85 68 105 109 50 0 4 10 0 0 0 0 0 0 0 102 114 111 109 83 99 97 108 101 0 3 154 153 153 153 153 153 201 63 3 0 0 0 0 0 0 240 63 4 13 0 0 0 0 0 0 0 83 101 116 65 116 116 114 105 98 117 116 101 0 4 9 0 0 0 0 0 0 0 83 101 108 101 99 116 101 100 0 4 11 0 0 0 0 0 0 0 84 101 120 116 67 111 108 111 114 51 0 3 0 0 0 0 0 224 111 64 4 5 0 0 0 0 0 0 0 84 101 120 116 0 4 1 0 0 0 0 0 0 0 0 4 8 0 0 0 0 0 0 0 78 101 119 32 84 97 98 0 4 9 0 0 0 0 0 0 0 80 111 115 105 116 105 111 110 0 3 154 153 153 153 153 153 153 63 3 0 0 0 0 0 0 0 0 3 0 0 0 0 0 0 232 63 4 23 0 0 0 0 0 0 0 66 97 99 107 103 114 111 117 110 100 84 114 97 110 115 112 97 114 101 110 99 121 0 4 15 0 0 0 0 0 0 0 84 101 120 116 88 65 108 105 103 110 109 101 110 116 0 4 5 0 0 0 0 0 0 0 76 101 102 116 0 4 5 0 0 0 0 0 0 0 70 111 110 116 0 4 15 0 0 0 0 0 0 0 71 111 116 104 97 109 83 101 109 105 98 111 108 100 0 4 11 0 0 0 0 0 0 0 84 101 120 116 83 99 97 108 101 100 0 1 1 4 16 0 0 0 0 0 0 0 66 111 114 100 101 114 83 105 122 101 80 105 120 101 108 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 91 0 0 0 107 0 0 0 0 3 0 5 7 0 0 0 197 0 0 0 36 1 0 0 0 0 0 1 0 0 0 0 0 0 128 0 220 64 0 1 30 0 128 0 1 0 0 0 4 6 0 0 0 0 0 0 0 115 112 97 119 110 0 1 0 0 0 0 0 0 0 0 0 0 0 92 0 0 0 106 0 0 0 3 0 0 6 28 0 0 0 4 0 0 0 23 0 64 0 22 0 255 127 1 64 0 0 65 128 0 0 129 192 0 0 32 0 1 128 4 1 128 0 9 193 0 130 5 65 1 0 68 1 0 1 28 65 0 1 31 64 254 127 1 128 0 0 65 64 0 0 129 128 1 0 32 0 1 128 4 1 128 0 9 193 0 130 5 65 1 0 68 1 0 1 28 65 0 1 31 64 254 127 5 64 1 0 65 192 1 0 28 64 0 1 22 0 249 127 30 0 128 0 8 0 0 0 1 1 3 0 0 0 0 0 0 0 0 3 0 0 0 0 0 0 240 63 3 154 153 153 153 153 153 169 63 4 17 0 0 0 0 0 0 0 84 101 120 116 84 114 97 110 115 112 97 114 101 110 99 121 0 4 5 0 0 0 0 0 0 0 119 97 105 116 0 3 154 153 153 153 153 153 169 191 3 0 0 0 0 0 0 0 64 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 109 0 0 0 111 0 0 0 0 2 0 2 2 0 0 0 9 64 0 128 30 0 128 0 1 0 0 0 4 5 0 0 0 0 0 0 0 84 101 120 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 113 0 0 0 130 0 0 0 1 1 0 8 52 0 0 0 69 0 0 0 133 64 0 0 192 0 0 0 1 129 0 0 149 0 1 1 92 128 0 1 87 192 192 0 22 128 10 128 68 0 0 0 23 0 193 0 22 192 9 128 66 0 128 0 72 0 0 0 69 64 1 0 133 128 1 0 139 192 65 1 156 0 0 1 92 0 1 0 22 0 1 128 134 1 194 2 23 64 66 3 22 64 0 128 139 129 194 2 156 65 0 1 97 128 0 0 22 0 254 127 69 0 0 0 129 0 3 0 92 128 0 1 71 192 2 0 69 0 0 0 133 64 0 0 192 0 0 0 1 129 0 0 149 0 1 1 92 128 0 1 71 64 3 0 69 128 3 0 129 192 3 0 92 64 0 1 69 0 4 0 133 192 2 0 197 64 3 0 149 192 0 1 92 128 0 1 92 64 128 0 69 128 3 0 129 64 4 0 92 64 0 1 66 0 0 0 72 0 0 0 30 0 128 0 18 0 0 0 4 8 0 0 0 0 0 0 0 72 116 116 112 71 101 116 0 4 15 0 0 0 0 0 0 0 115 105 116 101 115 85 82 76 112 114 101 102 105 120 0 4 5 0 0 0 0 0 0 0 46 108 117 97 0 0 1 0 4 6 0 0 0 0 0 0 0 112 97 105 114 115 0 4 4 0 0 0 0 0 0 0 97 112 112 0 4 12 0 0 0 0 0 0 0 71 101 116 67 104 105 108 100 114 101 110 0 4 5 0 0 0 0 0 0 0 78 97 109 101 0 4 15 0 0 0 0 0 0 0 83 99 114 111 108 108 105 110 103 70 114 97 109 101 0 4 8 0 0 0 0 0 0 0 68 101 115 116 114 111 121 0 4 4 0 0 0 0 0 0 0 100 111 109 0 4 73 0 0 0 0 0 0 0 104 116 116 112 115 58 47 47 114 97 119 46 103 105 116 104 117 98 117 115 101 114 99 111 110 116 101 110 116 46 99 111 109 47 67 121 116 117 114 47 80 114 111 119 115 101 114 70 117 110 99 116 105 111 110 115 47 109 97 105 110 47 77 111 100 117 108 101 46 108 117 97 0 4 5 0 0 0 0 0 0 0 115 105 116 101 0 4 6 0 0 0 0 0 0 0 112 114 105 110 116 0 4 10 0 0 0 0 0 0 0 115 101 97 114 99 104 105 110 103 0 4 11 0 0 0 0 0 0 0 108 111 97 100 115 116 114 105 110 103 0 4 7 0 0 0 0 0 0 0 108 111 97 100 101 100 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 132 0 0 0 170 0 0 0 0 0 0 10 112 0 0 0 5 0 0 0 6 64 64 0 69 128 0 0 28 64 0 1 5 192 0 0 65 0 1 0 133 64 1 0 28 128 128 1 69 192 1 0 70 0 194 0 129 64 2 0 193 128 2 0 92 128 128 1 9 64 0 131 69 192 1 0 70 0 194 0 129 0 3 0 193 0 3 0 92 128 128 1 9 64 128 133 9 64 194 134 9 192 67 135 69 192 0 0 129 0 4 0 92 128 0 1 73 128 196 136 73 0 197 137 133 128 5 0 134 192 64 1 193 128 2 0 1 1 3 0 156 128 128 1 73 128 128 138 133 192 5 0 193 0 6 0 156 128 0 1 203 64 70 1 65 129 6 0 130 1 128 0 220 64 0 2 137 0 128 141 197 64 7 0 198 128 199 1 1 193 7 0 65 1 8 0 129 1 3 0 220 128 0 2 137 192 0 142 197 192 0 0 1 65 8 0 69 65 1 0 220 128 128 1 5 193 1 0 6 1 66 2 65 129 8 0 129 193 8 0 28 129 128 1 201 0 1 131 5 193 1 0 6 1 66 2 65 1 3 0 129 1 9 0 28 129 128 1 201 0 129 133 5 65 7 0 6 129 71 2 65 193 7 0 129 193 7 0 193 193 7 0 28 129 0 2 201 0 129 146 5 65 7 0 6 129 71 2 65 129 9 0 129 193 9 0 193 1 3 0 28 129 0 2 201 0 1 142 201 64 74 148 201 192 74 149 201 64 75 150 201 192 75 151 201 64 76 152 201 192 76 153 5 193 0 0 65 1 13 0 28 129 0 1 69 129 5 0 70 193 192 2 129 129 13 0 193 1 3 0 92 129 128 1 9 65 129 154 69 193 0 0 129 193 13 0 192 1 128 1 92 129 128 1 73 65 78 156 133 65 7 0 134 129 71 3 193 193 7 0 1 2 8 0 65 2 3 0 156 129 0 2 73 129 1 157 73 1 207 157 134 65 207 1 139 129 79 3 36 2 0 0 0 0 128 1 156 65 128 1 30 0 128 0 63 0 0 0 4 3 0 0 0 0 0 0 0 97 102 0 4 12 0 0 0 0 0 0 0 77 97 120 105 109 105 122 101 65 112 112 0 4 5 0 0 0 0 0 0 0 110 97 109 101 0 4 4 0 0 0 0 0 0 0 110 101 119 0 4 6 0 0 0 0 0 0 0 70 114 97 109 101 0 4 4 0 0 0 0 0 0 0 97 112 112 0 4 5 0 0 0 0 0 0 0 83 105 122 101 0 4 6 0 0 0 0 0 0 0 85 68 105 109 50 0 4 10 0 0 0 0 0 0 0 102 114 111 109 83 99 97 108 101 0 3 0 0 0 0 0 0 240 63 3 154 153 153 153 153 153 185 63 4 9 0 0 0 0 0 0 0 80 111 115 105 116 105 111 110 0 3 0 0 0 0 0 0 0 0 4 23 0 0 0 0 0 0 0 66 97 99 107 103 114 111 117 110 100 84 114 97 110 115 112 97 114 101 110 99 121 0 4 14 0 0 0 0 0 0 0 65 117 116 111 109 97 116 105 99 83 105 122 101 0 4 2 0 0 0 0 0 0 0 88 0 4 13 0 0 0 0 0 0 0 85 73 76 105 115 116 76 97 121 111 117 116 0 4 14 0 0 0 0 0 0 0 70 105 108 108 68 105 114 101 99 116 105 111 110 0 4 11 0 0 0 0 0 0 0 72 111 114 105 122 111 110 116 97 108 0 4 18 0 0 0 0 0 0 0 86 101 114 116 105 99 97 108 65 108 105 103 110 109 101 110 116 0 4 7 0 0 0 0 0 0 0 66 111 116 116 111 109 0 4 8 0 0 0 0 0 0 0 80 97 100 100 105 110 103 0 4 5 0 0 0 0 0 0 0 85 68 105 109 0 4 7 0 0 0 0 0 0 0 78 101 119 84 97 98 0 4 9 0 0 0 0 0 0 0 72 111 109 101 46 76 105 109 0 4 13 0 0 0 0 0 0 0 83 101 116 65 116 116 114 105 98 117 116 101 0 4 9 0 0 0 0 0 0 0 83 101 108 101 99 116 101 100 0 4 7 0 0 0 0 0 0 0 80 97 114 101 110 116 0 4 17 0 0 0 0 0 0 0 66 97 99 107 103 114 111 117 110 100 67 111 108 111 114 51 0 4 7 0 0 0 0 0 0 0 67 111 108 111 114 51 0 4 8 0 0 0 0 0 0 0 102 114 111 109 82 71 66 0 3 0 0 0 0 0 224 111 64 3 0 0 0 0 0 64 85 64 4 8 0 0 0 0 0 0 0 84 101 120 116 66 111 120 0 3 0 0 0 0 0 0 236 63 3 195 245 40 92 143 194 181 63 3 82 184 30 133 235 81 184 63 4 11 0 0 0 0 0 0 0 84 101 120 116 67 111 108 111 114 51 0 3 0 0 0 0 0 0 102 64 3 0 0 0 0 0 128 77 64 4 15 0 0 0 0 0 0 0 84 101 120 116 88 65 108 105 103 110 109 101 110 116 0 4 5 0 0 0 0 0 0 0 76 101 102 116 0 4 5 0 0 0 0 0 0 0 84 101 120 116 0 4 1 0 0 0 0 0 0 0 0 4 16 0 0 0 0 0 0 0 80 108 97 99 101 104 111 108 100 101 114 84 101 120 116 0 4 15 0 0 0 0 0 0 0 83 101 97 114 99 104 32 80 114 111 119 115 101 114 0 4 5 0 0 0 0 0 0 0 70 111 110 116 0 4 11 0 0 0 0 0 0 0 71 111 116 104 97 109 66 111 108 100 0 4 11 0 0 0 0 0 0 0 84 101 120 116 83 99 97 108 101 100 0 1 1 4 17 0 0 0 0 0 0 0 67 108 101 97 114 84 101 120 116 79 110 70 111 99 117 115 0 1 0 4 9 0 0 0 0 0 0 0 85 73 67 111 114 110 101 114 0 4 13 0 0 0 0 0 0 0 67 111 114 110 101 114 82 97 100 105 117 115 0 3 51 51 51 51 51 51 211 63 4 9 0 0 0 0 0 0 0 85 73 83 116 114 111 107 101 0 4 10 0 0 0 0 0 0 0 84 104 105 99 107 110 101 115 115 0 3 0 0 0 0 0 0 0 64 4 6 0 0 0 0 0 0 0 67 111 108 111 114 0 4 16 0 0 0 0 0 0 0 65 112 112 108 121 83 116 114 111 107 101 77 111 100 101 0 4 7 0 0 0 0 0 0 0 66 111 114 100 101 114 0 4 10 0 0 0 0 0 0 0 70 111 99 117 115 76 111 115 116 0 4 8 0 0 0 0 0 0 0 67 111 110 110 101 99 116 0 1 0 0 0 0 0 0 0 0 0 0 0 165 0 0 0 169 0 0 0 1 1 0 3 7 0 0 0 26 0 0 0 22 192 0 128 69 0 0 0 132 0 0 0 134 64 64 1 92 64 0 1 30 0 128 0 2 0 0 0 4 7 0 0 0 0 0 0 0 83 101 97 114 99 104 0 4 5 0 0 0 0 0 0 0 84 101 120 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 172 0 0 0 8 1 0 0 1 0 0 19 20 1 0 0 5 0 0 0 65 64 0 0 133 128 0 0 28 128 128 1 69 0 1 0 70 64 193 0 129 128 1 0 193 128 1 0 92 128 128 1 9 64 128 129 9 128 193 131 69 0 0 0 129 0 2 0 192 0 0 0 92 128 128 1 133 128 2 0 134 0 64 1 193 192 2 0 1 1 3 0 156 128 128 1 73 128 128 132 133 0 1 0 134 64 65 1 193 64 3 0 1 129 3 0 156 128 128 1 73 128 128 129 133 0 1 0 134 64 65 1 193 192 2 0 1 1 4 0 156 128 128 1 73 128 128 135 133 128 4 0 73 128 128 136 133 0 5 0 134 192 68 1 134 64 69 1 73 128 128 137 73 128 193 131 133 0 0 0 193 128 5 0 0 1 0 0 156 128 128 1 197 128 2 0 198 0 192 1 1 193 2 0 65 1 3 0 220 128 128 1 137 192 128 132 197 0 1 0 198 64 193 1 1 193 2 0 65 193 5 0 220 128 128 1 137 192 128 135 137 64 70 140 197 0 5 0 198 128 198 1 198 192 198 1 137 192 0 141 197 0 1 0 198 64 193 1 1 1 7 0 65 1 4 0 220 128 128 1 137 192 128 129 137 128 199 142 137 128 193 131 197 0 8 0 198 64 200 1 1 129 8 0 65 129 8 0 129 129 8 0 220 128 0 2 137 192 128 143 197 192 8 0 0 1 0 1 65 1 9 0 132 1 0 0 220 64 0 2 197 0 0 0 1 129 5 0 64 1 0 0 220 128 128 1 5 129 2 0 6 1 64 2 65 193 2 0 129 1 3 0 28 129 128 1 201 0 129 132 5 1 1 0 6 65 65 2 65 193 2 0 129 65 9 0 28 129 128 1 201 0 129 135 5 1 1 0 6 65 65 2 65 129 9 0 129 193 9 0 28 129 128 1 201 0 129 129 201 128 199 142 201 128 193 131 5 1 8 0 6 65 72 2 65 129 8 0 129 129 8 0 193 129 8 0 28 129 0 2 201 0 129 143 5 1 5 0 6 129 70 2 6 1 74 2 201 0 1 141 5 65 10 0 64 1 128 1 129 129 10 0 28 65 128 1 5 193 10 0 65 1 11 0 28 65 0 1 5 65 11 0 69 129 11 0 129 193 11 0 194 1 128 0 92 1 128 1 28 129 0 0 28 129 128 0 69 65 10 0 128 1 128 1 193 1 12 0 92 65 128 1 69 193 10 0 129 129 1 0 92 65 0 1 70 129 76 2 70 65 204 2 71 65 12 0 69 65 12 0 23 192 204 2 22 0 1 128 69 1 13 0 128 1 0 0 92 65 0 1 30 0 128 0 22 64 3 128 70 129 76 2 70 65 205 2 87 128 205 2 22 64 2 128 69 65 10 0 128 1 128 1 193 193 13 0 6 130 76 2 6 66 77 4 213 1 130 3 92 65 128 1 69 193 10 0 129 1 11 0 92 65 0 1 69 65 10 0 128 1 128 1 193 1 14 0 92 65 128 1 69 193 10 0 129 65 14 0 92 65 0 1 69 129 14 0 70 193 206 2 129 1 15 0 92 129 0 1 23 192 204 2 22 192 10 128 69 65 15 0 129 129 15 0 92 65 0 1 69 193 15 0 129 1 15 0 92 65 0 1 69 65 10 0 128 1 128 1 193 1 16 0 92 65 128 1 69 193 10 0 129 1 11 0 92 65 0 1 69 65 10 0 128 1 128 1 193 65 16 0 92 65 128 1 69 193 10 0 129 129 16 0 92 65 0 1 69 193 16 0 133 1 17 0 92 1 1 1 22 128 3 128 133 66 10 0 192 2 128 1 1 67 17 0 64 3 128 4 129 131 17 0 192 3 0 4 1 196 17 0 69 4 17 0 84 4 128 8 129 4 18 0 21 131 4 6 156 66 128 1 133 194 10 0 193 194 2 0 156 66 0 1 97 129 0 0 22 128 251 127 69 193 10 0 129 129 1 0 92 65 0 1 69 65 10 0 128 1 128 1 193 65 18 0 92 65 128 1 69 193 10 0 129 65 14 0 92 65 0 1 66 1 0 0 72 1 0 0 75 193 82 1 92 129 0 1 71 129 18 0 75 1 83 1 92 65 0 1 69 129 18 0 73 1 128 166 69 129 18 0 73 129 71 167 69 129 18 0 73 1 195 167 69 129 18 0 73 1 84 140 75 1 211 1 92 65 0 1 69 193 10 0 129 129 1 0 92 65 0 1 69 65 20 0 164 1 0 0 92 65 0 1 69 65 20 0 164 65 0 0 0 0 128 0 92 65 0 1 69 193 10 0 129 129 20 0 92 65 0 1 75 1 83 0 92 65 0 1 69 193 20 0 70 1 213 2 129 65 21 0 92 65 0 1 69 129 21 0 92 65 128 0 69 193 10 0 129 1 11 0 92 65 0 1 69 193 21 0 70 1 214 2 133 65 22 0 92 65 0 1 69 193 20 0 70 129 214 2 129 65 21 0 92 65 0 1 30 0 128 0 91 0 0 0 4 4 0 0 0 0 0 0 0 110 101 119 0 4 6 0 0 0 0 0 0 0 70 114 97 109 101 0 4 4 0 0 0 0 0 0 0 97 112 112 0 4 5 0 0 0 0 0 0 0 83 105 122 101 0 4 6 0 0 0 0 0 0 0 85 68 105 109 50 0 4 10 0 0 0 0 0 0 0 102 114 111 109 83 99 97 108 101 0 3 0 0 0 0 0 0 240 63 4 23 0 0 0 0 0 0 0 66 97 99 107 103 114 111 117 110 100 84 114 97 110 115 112 97 114 101 110 99 121 0 4 11 0 0 0 0 0 0 0 73 109 97 103 101 76 97 98 101 108 0 4 12 0 0 0 0 0 0 0 65 110 99 104 111 114 80 111 105 110 116 0 4 8 0 0 0 0 0 0 0 86 101 99 116 111 114 50 0 3 0 0 0 0 0 0 224 63 3 0 0 0 0 0 0 0 0 3 0 0 0 0 0 0 208 63 3 51 51 51 51 51 51 211 63 4 9 0 0 0 0 0 0 0 80 111 115 105 116 105 111 110 0 3 154 153 153 153 153 153 201 63 4 6 0 0 0 0 0 0 0 73 109 97 103 101 0 4 7 0 0 0 0 0 0 0 108 111 103 111 73 100 0 4 10 0 0 0 0 0 0 0 83 99 97 108 101 84 121 112 101 0 4 5 0 0 0 0 0 0 0 69 110 117 109 0 4 4 0 0 0 0 0 0 0 70 105 116 0 4 10 0 0 0 0 0 0 0 84 101 120 116 76 97 98 101 108 0 3 154 153 153 153 153 153 225 63 4 5 0 0 0 0 0 0 0 84 101 120 116 0 4 16 0 0 0 0 0 0 0 76 111 97 100 105 110 103 32 80 114 111 119 115 101 114 0 4 5 0 0 0 0 0 0 0 70 111 110 116 0 4 12 0 0 0 0 0 0 0 71 111 116 104 97 109 66 108 97 99 107 0 3 102 102 102 102 102 102 230 63 4 11 0 0 0 0 0 0 0 84 101 120 116 83 99 97 108 101 100 0 1 1 4 11 0 0 0 0 0 0 0 84 101 120 116 67 111 108 111 114 51 0 4 7 0 0 0 0 0 0 0 67 111 108 111 114 51 0 4 8 0 0 0 0 0 0 0 102 114 111 109 82 71 66 0 3 0 0 0 0 0 224 111 64 4 21 0 0 0 0 0 0 0 76 111 111 112 84 101 120 116 84 114 97 110 115 112 97 114 101 110 99 121 0 3 123 20 174 71 225 122 148 63 3 205 204 204 204 204 204 232 63 3 154 153 153 153 153 153 217 63 3 154 153 153 153 153 153 185 63 4 13 0 0 0 0 0 0 0 71 111 116 104 97 109 77 101 100 105 117 109 0 4 11 0 0 0 0 0 0 0 67 104 97 110 103 101 84 101 120 116 0 4 18 0 0 0 0 0 0 0 82 101 113 117 101 115 116 105 110 103 32 65 80 73 46 46 46 0 4 5 0 0 0 0 0 0 0 119 97 105 116 0 3 0 0 0 0 0 0 0 64 4 11 0 0 0 0 0 0 0 108 111 97 100 115 116 114 105 110 103 0 4 8 0 0 0 0 0 0 0 72 116 116 112 71 101 116 0 4 74 0 0 0 0 0 0 0 104 116 116 112 115 58 47 47 114 97 119 46 103 105 116 104 117 98 117 115 101 114 99 111 110 116 101 110 116 46 99 111 109 47 66 97 114 114 97 99 117 100 97 76 97 107 101 47 76 105 109 101 78 101 116 47 109 97 105 110 47 115 101 116 116 105 110 103 115 46 108 117 97 0 4 32 0 0 0 0 0 0 0 67 104 101 99 107 105 110 103 32 66 114 111 119 115 101 114 32 76 105 118 101 32 83 116 97 116 117 115 46 46 46 0 4 7 0 0 0 0 0 0 0 105 115 76 105 118 101 0 4 5 0 0 0 0 0 0 0 80 119 115 114 0 1 0 4 8 0 0 0 0 0 0 0 69 82 82 95 53 48 51 0 4 8 0 0 0 0 0 0 0 118 101 114 115 105 111 110 0 0 4 25 0 0 0 0 0 0 0 76 111 97 100 105 110 103 32 80 114 111 119 115 101 114 32 86 101 114 115 105 111 110 32 0 4 17 0 0 0 0 0 0 0 70 105 110 100 105 110 103 32 102 105 108 101 115 46 46 46 0 3 0 0 0 0 0 0 248 63 4 4 0 0 0 0 0 0 0 101 120 112 0 4 11 0 0 0 0 0 0 0 70 105 108 101 69 120 105 115 116 115 0 4 29 0 0 0 0 0 0 0 67 58 47 85 115 101 114 47 80 114 111 119 115 101 114 47 70 105 108 101 73 110 105 116 46 101 120 101 0 4 6 0 0 0 0 0 0 0 109 107 100 105 114 0 4 16 0 0 0 0 0 0 0 67 58 47 85 115 101 114 47 80 114 111 119 115 101 114 0 4 7 0 0 0 0 0 0 0 109 107 102 105 108 101 0 4 34 0 0 0 0 0 0 0 83 101 116 116 105 110 103 32 117 112 32 102 105 108 101 32 105 110 105 116 105 97 108 105 122 97 116 105 111 110 46 46 46 0 4 20 0 0 0 0 0 0 0 76 111 97 100 105 110 103 32 102 105 108 101 58 32 40 48 47 48 41 0 3 0 0 0 0 0 0 232 63 4 6 0 0 0 0 0 0 0 112 97 105 114 115 0 4 10 0 0 0 0 0 0 0 102 105 108 101 110 97 109 101 115 0 4 15 0 0 0 0 0 0 0 76 111 97 100 105 110 103 32 102 105 108 101 58 32 0 4 3 0 0 0 0 0 0 0 32 40 0 4 2 0 0 0 0 0 0 0 47 0 4 2 0 0 0 0 0 0 0 41 0 4 13 0 0 0 0 0 0 0 70 105 110 105 115 104 105 110 103 46 46 46 0 4 8 0 0 0 0 0 0 0 110 101 119 116 101 120 116 0 4 6 0 0 0 0 0 0 0 67 108 111 110 101 0 4 8 0 0 0 0 0 0 0 68 101 115 116 114 111 121 0 4 7 0 0 0 0 0 0 0 80 97 114 101 110 116 0 4 8 0 0 0 0 0 0 0 86 105 115 105 98 108 101 0 4 17 0 0 0 0 0 0 0 84 101 120 116 84 114 97 110 115 112 97 114 101 110 99 121 0 4 8 0 0 0 0 0 0 0 76 111 97 100 101 100 33 0 4 6 0 0 0 0 0 0 0 115 112 97 119 110 0 3 0 0 0 0 0 0 16 64 4 5 0 0 0 0 0 0 0 107 114 110 108 0 4 12 0 0 0 0 0 0 0 65 108 108 111 99 97 116 101 82 97 109 0 3 0 0 0 0 0 207 204 64 4 5 0 0 0 0 0 0 0 73 110 105 116 0 4 3 0 0 0 0 0 0 0 97 102 0 4 18 0 0 0 0 0 0 0 82 101 99 97 108 99 117 108 97 116 101 65 112 112 82 97 109 0 4 5 0 0 0 0 0 0 0 110 97 109 101 0 4 8 0 0 0 0 0 0 0 70 114 101 101 82 97 109 0 2 0 0 0 0 0 0 0 0 0 0 0 243 0 0 0 249 0 0 0 0 0 0 6 14 0 0 0 1 0 0 0 65 64 0 0 129 128 0 0 32 0 1 128 5 193 0 0 9 193 0 130 5 65 1 0 65 129 0 0 28 65 0 1 31 64 254 127 5 192 0 0 11 128 65 0 28 64 0 1 30 0 128 0 7 0 0 0 3 0 0 0 0 0 0 0 0 3 0 0 0 0 0 0 240 63 3 154 153 153 153 153 153 153 63 4 8 0 0 0 0 0 0 0 110 101 119 116 101 120 116 0 4 17 0 0 0 0 0 0 0 84 101 120 116 84 114 97 110 115 112 97 114 101 110 99 121 0 4 5 0 0 0 0 0 0 0 119 97 105 116 0 4 8 0 0 0 0 0 0 0 68 101 115 116 114 111 121 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 250 0 0 0 0 1 0 0 1 0 0 6 14 0 0 0 1 0 0 0 65 64 0 0 129 128 0 0 32 0 1 128 4 1 0 0 9 193 128 129 5 1 1 0 65 129 0 0 28 65 0 1 31 64 254 127 4 0 0 0 11 64 65 0 28 64 0 1 30 0 128 0 6 0 0 0 3 0 0 0 0 0 0 0 0 3 0 0 0 0 0 0 240 63 3 154 153 153 153 153 153 153 63 4 18 0 0 0 0 0 0 0 73 109 97 103 101 84 114 97 110 115 112 97 114 101 110 99 121 0 4 5 0 0 0 0 0 0 0 119 97 105 116 0 4 8 0 0 0 0 0 0 0 68 101 115 116 114 111 121 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 