76 69 70 0 0 0 0 0 1 0 0 0 0 0 0 0 57 66 105 116 66 121 116 101 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 97 57 57 51 50 102 52 53 102 48 51 97 100 52 57 55 54 51 57 51 48 50 98 53 48 51 50 51 53 56 50 56 52 51 55 55 53 51 51 56 97 97 97 55 53 98 55 50 48 49 97 55 99 98 97 100 52 50 57 52 97 55 48 57 27 76 117 97 81 0 1 4 8 4 8 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 2 12 194 0 0 0 5 0 0 0 65 64 0 0 28 128 0 1 65 128 0 0 129 192 0 0 193 0 1 0 5 65 1 0 65 129 1 0 128 1 0 0 28 129 128 1 9 1 194 131 69 129 2 0 70 193 194 2 129 1 3 0 193 65 3 0 92 129 128 1 9 65 129 132 69 129 2 0 70 193 194 2 129 193 3 0 193 1 4 0 92 129 128 1 9 65 1 135 9 129 196 136 9 1 197 137 9 129 197 138 69 1 6 0 70 65 198 2 129 129 6 0 193 129 6 0 1 130 6 0 92 129 0 2 9 65 129 139 69 1 6 0 70 65 198 2 129 129 6 0 193 129 6 0 1 130 6 0 92 129 0 2 9 65 129 141 69 1 6 0 70 65 198 2 129 65 7 0 193 65 7 0 1 66 7 0 92 129 0 2 9 65 1 142 69 65 1 0 129 129 1 0 192 1 0 0 92 129 128 1 73 129 199 131 133 129 2 0 134 193 66 3 193 1 3 0 1 66 3 0 156 129 128 1 73 129 129 132 133 129 2 0 134 193 66 3 193 193 3 0 1 194 7 0 156 129 128 1 73 129 1 135 73 1 200 136 73 1 197 137 73 129 197 138 133 1 6 0 134 65 70 3 193 129 6 0 1 130 6 0 65 130 6 0 156 129 0 2 73 129 129 139 133 1 6 0 134 65 70 3 193 129 6 0 1 130 6 0 65 130 6 0 156 129 0 2 73 129 129 141 133 1 6 0 134 65 70 3 193 65 7 0 1 66 7 0 65 66 7 0 156 129 0 2 73 129 1 142 133 65 1 0 193 65 8 0 0 2 0 0 156 129 128 1 137 129 200 131 197 129 2 0 198 193 194 3 1 194 3 0 65 66 3 0 220 129 128 1 137 193 129 132 197 129 2 0 198 193 194 3 1 194 8 0 65 66 3 0 220 129 128 1 137 193 1 135 193 1 9 0 0 2 128 0 213 1 130 3 137 193 129 136 137 1 197 137 137 129 197 138 197 1 6 0 198 65 198 3 1 130 6 0 65 130 6 0 129 130 6 0 220 129 0 2 137 193 129 139 197 1 6 0 198 65 198 3 1 130 6 0 65 130 6 0 129 130 6 0 220 129 0 2 137 193 129 141 197 1 6 0 198 65 198 3 1 66 7 0 65 66 7 0 129 66 7 0 220 129 0 2 137 193 1 142 197 65 1 0 1 66 8 0 64 2 0 0 220 129 128 1 201 65 201 131 5 130 2 0 6 194 66 4 65 194 8 0 129 66 3 0 28 130 128 1 201 1 130 132 5 130 2 0 6 194 66 4 65 130 9 0 129 194 9 0 28 130 128 1 201 1 2 135 1 2 10 0 64 2 0 1 21 66 2 4 201 1 130 136 201 1 197 137 201 129 197 138 5 2 6 0 6 66 70 4 65 130 6 0 129 130 6 0 193 130 6 0 28 130 0 2 201 1 130 139 5 2 6 0 6 66 70 4 65 130 6 0 129 130 6 0 193 130 6 0 28 130 0 2 201 1 130 141 5 2 6 0 6 66 70 4 65 66 7 0 129 66 7 0 193 66 7 0 28 130 0 2 201 1 2 142 6 66 74 2 11 130 74 4 164 2 0 0 0 0 128 0 0 0 0 1 0 0 0 3 28 66 128 1 6 66 202 2 11 130 74 4 164 66 0 0 0 0 128 0 0 0 128 1 0 0 0 1 0 0 128 3 0 0 0 3 0 0 128 2 28 66 128 1 30 0 128 0 43 0 0 0 4 10 0 0 0 0 0 0 0 99 114 101 97 116 101 97 112 112 0 4 13 0 0 0 0 0 0 0 67 108 105 99 107 101 114 32 71 97 109 101 0 3 0 0 0 0 0 0 0 0 3 0 0 0 0 0 0 240 63 3 0 0 0 0 0 0 0 64 4 4 0 0 0 0 0 0 0 110 101 119 0 4 11 0 0 0 0 0 0 0 84 101 120 116 66 117 116 116 111 110 0 4 5 0 0 0 0 0 0 0 78 97 109 101 0 4 11 0 0 0 0 0 0 0 77 97 105 110 66 117 116 116 111 110 0 4 5 0 0 0 0 0 0 0 83 105 122 101 0 4 6 0 0 0 0 0 0 0 85 68 105 109 50 0 4 10 0 0 0 0 0 0 0 102 114 111 109 83 99 97 108 101 0 3 154 153 153 153 153 153 217 63 3 154 153 153 153 153 153 185 63 4 9 0 0 0 0 0 0 0 80 111 115 105 116 105 111 110 0 3 51 51 51 51 51 51 211 63 3 0 0 0 0 0 0 224 63 4 5 0 0 0 0 0 0 0 84 101 120 116 0 4 10 0 0 0 0 0 0 0 67 108 105 99 107 32 77 101 33 0 4 11 0 0 0 0 0 0 0 84 101 120 116 83 99 97 108 101 100 0 1 1 4 5 0 0 0 0 0 0 0 70 111 110 116 0 4 7 0 0 0 0 0 0 0 71 111 116 104 97 109 0 4 17 0 0 0 0 0 0 0 66 97 99 107 103 114 111 117 110 100 67 111 108 111 114 51 0 4 7 0 0 0 0 0 0 0 67 111 108 111 114 51 0 4 8 0 0 0 0 0 0 0 102 114 111 109 82 71 66 0 3 0 0 0 0 0 128 70 64 4 13 0 0 0 0 0 0 0 66 111 114 100 101 114 67 111 108 111 114 51 0 4 11 0 0 0 0 0 0 0 84 101 120 116 67 111 108 111 114 51 0 3 0 0 0 0 0 224 111 64 4 14 0 0 0 0 0 0 0 85 112 103 114 97 100 101 66 117 116 116 111 110 0 3 102 102 102 102 102 102 230 63 4 19 0 0 0 0 0 0 0 85 112 103 114 97 100 101 32 77 117 108 116 105 112 108 105 101 114 0 4 10 0 0 0 0 0 0 0 84 101 120 116 76 97 98 101 108 0 4 7 0 0 0 0 0 0 0 67 108 105 99 107 115 0 3 102 102 102 102 102 102 214 63 4 9 0 0 0 0 0 0 0 67 108 105 99 107 115 58 32 0 4 4 0 0 0 0 0 0 0 77 85 76 0 3 205 204 204 204 204 204 212 63 3 205 204 204 204 204 204 204 63 4 16 0 0 0 0 0 0 0 77 117 108 116 105 112 108 105 99 97 116 111 114 58 32 0 4 18 0 0 0 0 0 0 0 77 111 117 115 101 66 117 116 116 111 110 49 67 108 105 99 107 0 4 8 0 0 0 0 0 0 0 67 111 110 110 101 99 116 0 2 0 0 0 0 0 0 0 0 0 0 0 55 0 0 0 58 0 0 0 3 0 0 3 11 0 0 0 4 0 0 0 68 0 128 0 78 64 0 128 12 64 0 0 8 0 0 0 4 0 0 1 65 128 0 0 132 0 0 0 85 128 128 0 9 64 128 128 30 0 128 0 3 0 0 0 3 0 0 0 0 0 0 240 63 4 5 0 0 0 0 0 0 0 84 101 120 116 0 4 9 0 0 0 0 0 0 0 67 108 105 99 107 115 58 32 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 60 0 0 0 73 0 0 0 6 0 0 4 44 0 0 0 4 0 0 0 68 0 128 0 25 0 128 0 22 192 5 128 4 0 0 0 68 0 128 0 13 64 0 0 8 0 0 0 4 0 0 1 8 0 128 0 4 0 0 1 14 0 64 0 69 64 0 0 70 128 192 0 140 192 64 0 92 128 0 1 72 0 0 1 68 0 128 1 129 64 1 0 196 0 0 1 149 192 0 1 73 128 0 130 68 0 0 2 129 128 1 0 196 0 0 0 149 192 0 1 73 128 0 130 22 128 3 128 4 0 0 0 68 0 128 0 24 64 0 0 22 128 2 128 4 0 128 2 65 192 1 0 132 0 128 0 193 0 2 0 85 192 128 0 9 64 0 130 5 64 2 0 65 128 2 0 28 64 0 1 4 0 128 2 9 192 66 130 30 0 128 0 12 0 0 0 3 47 221 36 6 129 149 4 64 4 5 0 0 0 0 0 0 0 109 97 116 104 0 4 6 0 0 0 0 0 0 0 102 108 111 111 114 0 3 0 0 0 0 0 0 240 63 4 5 0 0 0 0 0 0 0 84 101 120 116 0 4 16 0 0 0 0 0 0 0 77 117 108 116 105 112 108 105 99 97 116 111 114 58 32 0 4 9 0 0 0 0 0 0 0 67 108 105 99 107 115 58 32 0 4 10 0 0 0 0 0 0 0 89 111 117 32 110 101 101 100 32 0 4 9 0 0 0 0 0 0 0 32 67 108 105 99 107 115 33 0 4 5 0 0 0 0 0 0 0 119 97 105 116 0 3 0 0 0 0 0 0 0 64 4 19 0 0 0 0 0 0 0 85 112 103 114 97 100 101 32 77 117 108 116 105 112 108 105 101 114 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 