76 69 70 0 0 0 0 0 1 0 0 0 0 0 0 0 57 66 105 116 66 121 116 101 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 52 101 52 53 100 102 56 102 57 48 51 49 51 101 48 100 55 100 97 54 55 56 53 53 101 52 98 50 52 99 56 101 54 97 57 56 55 49 54 49 54 98 56 98 51 52 51 52 48 57 52 98 48 101 55 98 53 98 49 102 100 52 55 48 27 76 117 97 81 0 1 4 8 4 8 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 2 9 92 0 0 0 10 0 0 0 69 0 0 0 70 64 192 0 129 128 0 0 92 128 0 1 133 0 0 0 134 192 64 1 192 0 128 0 1 1 1 0 156 128 128 1 137 128 193 130 197 0 2 0 198 64 194 1 1 129 2 0 65 193 2 0 220 128 128 1 137 192 128 131 197 64 3 0 198 128 195 1 1 193 3 0 65 1 4 0 129 1 4 0 220 128 0 2 137 192 0 134 137 128 196 136 197 192 4 0 1 1 5 0 220 64 0 1 197 0 0 0 198 192 192 1 0 1 128 0 65 65 5 0 220 128 128 1 201 128 193 130 201 128 197 136 5 1 2 0 6 65 66 2 65 193 5 0 129 1 6 0 28 129 128 1 201 0 129 131 5 65 3 0 6 129 67 2 65 193 3 0 129 1 4 0 193 1 4 0 28 129 0 2 201 0 1 134 5 1 2 0 6 65 66 2 65 1 4 0 129 193 2 0 28 129 128 1 201 0 129 140 6 129 198 1 11 193 70 2 164 1 0 0 0 0 128 0 28 65 128 1 5 1 0 0 6 193 64 2 64 1 128 0 129 65 5 0 28 129 128 1 9 129 193 130 9 1 199 136 69 1 2 0 70 65 194 2 129 193 5 0 193 1 6 0 92 129 128 1 9 65 129 131 69 65 3 0 70 129 195 2 129 1 4 0 193 193 3 0 1 2 4 0 92 129 0 2 9 65 1 134 69 1 2 0 70 65 194 2 129 193 5 0 193 193 2 0 92 129 128 1 9 65 129 140 70 129 70 2 75 193 198 2 228 65 0 0 0 0 128 0 0 0 0 0 92 65 128 1 30 0 128 0 29 0 0 0 4 5 0 0 0 0 0 0 0 76 105 109 101 0 4 13 0 0 0 0 0 0 0 67 114 101 97 116 101 87 105 110 100 111 119 0 4 12 0 0 0 0 0 0 0 68 105 115 99 108 97 105 109 101 114 33 0 4 9 0 0 0 0 0 0 0 67 114 101 97 116 101 85 73 0 4 10 0 0 0 0 0 0 0 84 101 120 116 76 97 98 101 108 0 4 11 0 0 0 0 0 0 0 84 101 120 116 83 99 97 108 101 100 0 1 1 4 5 0 0 0 0 0 0 0 83 105 122 101 0 4 6 0 0 0 0 0 0 0 85 68 105 109 50 0 4 10 0 0 0 0 0 0 0 102 114 111 109 83 99 97 108 101 0 3 0 0 0 0 0 0 240 63 3 205 204 204 204 204 204 236 63 4 17 0 0 0 0 0 0 0 66 97 99 107 103 114 111 117 110 100 67 111 108 111 114 51 0 4 7 0 0 0 0 0 0 0 67 111 108 111 114 51 0 4 8 0 0 0 0 0 0 0 102 114 111 109 82 71 66 0 3 0 0 0 0 0 224 111 64 3 0 0 0 0 0 0 0 0 4 5 0 0 0 0 0 0 0 84 101 120 116 0 4 97 0 0 0 0 0 0 0 68 73 83 67 76 65 73 77 69 82 33 32 66 121 32 99 111 110 116 105 110 117 105 110 103 32 32 121 111 117 32 117 110 100 101 114 115 116 97 110 100 32 116 104 97 116 32 97 116 32 97 110 121 32 116 105 109 101 32 97 108 108 32 111 102 32 121 111 117 114 32 119 105 110 100 111 119 115 32 99 111 117 108 100 32 98 101 32 99 108 101 97 114 101 100 46 0 4 5 0 0 0 0 0 0 0 119 97 105 116 0 3 0 0 0 0 0 0 32 64 4 11 0 0 0 0 0 0 0 84 101 120 116 66 117 116 116 111 110 0 4 27 0 0 0 0 0 0 0 73 32 100 111 32 110 111 116 32 119 105 115 104 32 116 111 32 99 111 110 116 105 110 117 101 46 0 3 0 0 0 0 0 0 224 63 3 154 153 153 153 153 153 185 63 4 9 0 0 0 0 0 0 0 80 111 115 105 116 105 111 110 0 4 18 0 0 0 0 0 0 0 77 111 117 115 101 66 117 116 116 111 110 49 67 108 105 99 107 0 4 8 0 0 0 0 0 0 0 67 111 110 110 101 99 116 0 4 20 0 0 0 0 0 0 0 73 32 119 105 115 104 32 116 111 32 99 111 110 116 105 110 117 101 46 0 2 0 0 0 0 0 0 0 0 0 0 0 16 0 0 0 18 0 0 0 1 1 0 3 10 0 0 0 69 0 0 0 129 64 0 0 92 128 0 1 70 128 192 0 132 0 0 0 134 192 64 1 134 0 65 1 134 0 65 1 92 64 0 1 30 0 128 0 5 0 0 0 4 8 0 0 0 0 0 0 0 108 111 97 100 108 105 98 0 4 19 0 0 0 0 0 0 0 65 112 112 108 105 99 97 116 105 111 110 72 97 110 100 108 101 114 0 4 12 0 0 0 0 0 0 0 69 120 105 116 80 114 111 99 101 115 115 0 4 7 0 0 0 0 0 0 0 80 97 114 101 110 116 0 4 6 0 0 0 0 0 0 0 86 97 108 117 101 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 26 0 0 0 95 2 0 0 2 1 0 10 101 0 0 0 69 0 0 0 129 64 0 0 92 128 0 1 70 128 192 0 132 0 0 0 134 192 64 1 134 0 65 1 134 0 65 1 92 64 0 1 66 0 128 0 133 64 1 0 134 128 65 1 193 192 1 0 156 128 0 1 197 64 1 0 198 0 194 1 0 1 0 1 65 65 2 0 220 128 128 1 201 192 66 133 5 65 3 0 6 129 67 2 65 193 3 0 129 1 4 0 28 129 128 1 201 0 1 134 5 129 4 0 6 193 68 2 65 1 5 0 129 65 5 0 193 65 5 0 28 129 0 2 201 0 129 136 201 192 69 139 5 1 6 0 65 65 6 0 28 65 0 1 5 65 1 0 6 1 66 2 64 1 0 1 129 129 6 0 28 129 128 1 9 193 66 133 9 193 70 139 69 65 3 0 70 129 195 2 129 1 7 0 193 65 7 0 92 129 128 1 9 65 1 134 69 129 4 0 70 193 196 2 129 1 5 0 193 65 5 0 1 66 5 0 92 129 0 2 9 65 129 136 69 65 3 0 70 129 195 2 129 65 5 0 193 1 4 0 92 129 128 1 9 65 1 143 70 193 71 2 75 1 200 2 228 1 0 0 0 0 0 1 92 65 128 1 69 65 1 0 70 1 194 2 128 1 0 1 193 129 6 0 92 129 128 1 73 193 66 133 73 65 72 139 133 65 3 0 134 129 67 3 193 1 7 0 1 66 7 0 156 129 128 1 73 129 1 134 133 129 4 0 134 193 68 3 193 65 5 0 1 2 5 0 65 66 5 0 156 129 0 2 73 129 129 136 133 65 3 0 134 129 67 3 193 1 7 0 1 2 4 0 156 129 128 1 73 129 1 143 134 193 199 2 139 1 72 3 36 66 0 0 0 0 0 1 4 0 128 0 156 65 128 1 30 0 128 0 34 0 0 0 4 8 0 0 0 0 0 0 0 108 111 97 100 108 105 98 0 4 19 0 0 0 0 0 0 0 65 112 112 108 105 99 97 116 105 111 110 72 97 110 100 108 101 114 0 4 12 0 0 0 0 0 0 0 69 120 105 116 80 114 111 99 101 115 115 0 4 7 0 0 0 0 0 0 0 80 97 114 101 110 116 0 4 6 0 0 0 0 0 0 0 86 97 108 117 101 0 4 5 0 0 0 0 0 0 0 76 105 109 101 0 4 13 0 0 0 0 0 0 0 67 114 101 97 116 101 87 105 110 100 111 119 0 4 14 0 0 0 0 0 0 0 68 105 115 99 108 97 105 109 101 114 32 50 33 0 4 9 0 0 0 0 0 0 0 67 114 101 97 116 101 85 73 0 4 10 0 0 0 0 0 0 0 84 101 120 116 76 97 98 101 108 0 4 11 0 0 0 0 0 0 0 84 101 120 116 83 99 97 108 101 100 0 1 1 4 5 0 0 0 0 0 0 0 83 105 122 101 0 4 6 0 0 0 0 0 0 0 85 68 105 109 50 0 4 10 0 0 0 0 0 0 0 102 114 111 109 83 99 97 108 101 0 3 0 0 0 0 0 0 240 63 3 205 204 204 204 204 204 236 63 4 17 0 0 0 0 0 0 0 66 97 99 107 103 114 111 117 110 100 67 111 108 111 114 51 0 4 7 0 0 0 0 0 0 0 67 111 108 111 114 51 0 4 8 0 0 0 0 0 0 0 102 114 111 109 82 71 66 0 3 0 0 0 0 0 224 111 64 3 0 0 0 0 0 0 0 0 4 5 0 0 0 0 0 0 0 84 101 120 116 0 4 142 0 0 0 0 0 0 0 68 73 83 67 76 65 73 77 69 82 33 32 66 121 32 99 111 110 116 105 110 117 105 110 103 32 32 121 111 117 32 117 110 100 101 114 115 116 97 110 100 32 116 104 97 116 32 97 116 32 97 110 121 32 116 105 109 101 32 121 111 117 32 109 97 121 32 110 111 116 32 98 101 32 97 98 108 101 32 116 111 32 100 111 32 97 110 121 116 104 105 110 103 32 102 111 114 32 116 101 109 112 111 114 97 114 105 97 108 32 97 109 111 117 110 116 115 32 111 102 32 116 105 109 101 32 119 105 116 104 32 110 111 32 101 115 99 97 112 101 46 0 4 5 0 0 0 0 0 0 0 119 97 105 116 0 3 0 0 0 0 0 0 32 64 4 11 0 0 0 0 0 0 0 84 101 120 116 66 117 116 116 111 110 0 4 27 0 0 0 0 0 0 0 73 32 100 111 32 110 111 116 32 119 105 115 104 32 116 111 32 99 111 110 116 105 110 117 101 46 0 3 0 0 0 0 0 0 224 63 3 154 153 153 153 153 153 185 63 4 9 0 0 0 0 0 0 0 80 111 115 105 116 105 111 110 0 4 18 0 0 0 0 0 0 0 77 111 117 115 101 66 117 116 116 111 110 49 67 108 105 99 107 0 4 8 0 0 0 0 0 0 0 67 111 110 110 101 99 116 0 4 20 0 0 0 0 0 0 0 73 32 119 105 115 104 32 116 111 32 99 111 110 116 105 110 117 101 46 0 2 0 0 0 0 0 0 0 0 0 0 0 43 0 0 0 45 0 0 0 1 1 0 3 10 0 0 0 69 0 0 0 129 64 0 0 92 128 0 1 70 128 192 0 132 0 0 0 134 192 64 1 134 0 65 1 134 0 65 1 92 64 0 1 30 0 128 0 5 0 0 0 4 8 0 0 0 0 0 0 0 108 111 97 100 108 105 98 0 4 19 0 0 0 0 0 0 0 65 112 112 108 105 99 97 116 105 111 110 72 97 110 100 108 101 114 0 4 12 0 0 0 0 0 0 0 69 120 105 116 80 114 111 99 101 115 115 0 4 7 0 0 0 0 0 0 0 80 97 114 101 110 116 0 4 6 0 0 0 0 0 0 0 86 97 108 117 101 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 53 0 0 0 94 2 0 0 2 1 0 25 225 0 0 0 69 0 0 0 129 64 0 0 92 128 0 1 70 128 192 0 132 0 0 0 134 192 64 1 134 0 65 1 134 0 65 1 92 64 0 1 66 0 0 0 133 64 1 0 134 128 65 1 193 192 1 0 1 1 2 0 156 128 128 1 202 0 128 5 1 65 2 0 65 129 2 0 129 193 2 0 193 1 3 0 1 66 3 0 65 130 3 0 129 194 3 0 193 2 4 0 1 67 4 0 65 131 4 0 129 195 4 0 226 64 128 5 10 1 128 5 65 1 5 0 129 65 5 0 193 1 5 0 1 2 5 0 65 66 5 0 129 2 5 0 193 2 5 0 1 3 5 0 65 67 5 0 129 67 5 0 193 3 5 0 34 65 128 5 65 129 5 0 130 1 0 0 228 1 0 0 5 194 5 0 65 2 6 0 28 66 0 1 36 66 0 0 69 194 5 0 129 66 6 0 92 66 0 1 69 66 1 0 70 130 198 4 128 2 0 1 193 194 6 0 92 130 128 1 133 66 7 0 134 130 71 5 193 194 7 0 1 3 8 0 65 67 8 0 129 3 8 0 156 130 128 2 73 130 2 142 133 66 7 0 134 130 71 5 193 2 8 0 1 3 8 0 65 195 8 0 129 3 8 0 156 130 128 2 73 130 2 145 73 66 73 146 133 194 9 0 134 2 74 5 193 66 10 0 1 131 10 0 65 3 8 0 156 130 0 2 73 130 2 147 73 2 203 149 133 194 9 0 134 2 74 5 193 130 10 0 1 131 10 0 65 131 10 0 156 130 0 2 73 130 130 150 73 194 75 151 133 66 1 0 134 130 70 5 192 2 0 1 1 195 6 0 156 130 128 1 197 66 7 0 198 130 199 5 1 195 7 0 65 3 8 0 129 67 8 0 193 3 8 0 220 130 128 2 137 194 2 142 137 2 76 146 197 194 9 0 198 2 202 5 1 131 10 0 65 3 8 0 129 3 8 0 220 130 0 2 137 194 2 147 197 66 7 0 198 130 199 5 1 67 12 0 65 3 8 0 129 195 8 0 193 3 8 0 220 130 128 2 137 194 2 145 137 2 203 149 197 194 9 0 198 2 202 5 1 131 10 0 65 131 10 0 129 131 10 0 220 130 0 2 137 194 130 150 137 130 76 151 197 66 1 0 198 130 198 5 0 3 0 1 65 195 12 0 220 130 128 1 5 67 7 0 6 131 71 6 65 131 5 0 129 3 8 0 193 67 8 0 1 4 8 0 28 131 128 2 201 2 3 142 5 67 7 0 6 131 71 6 65 3 8 0 129 3 8 0 193 3 8 0 1 4 8 0 28 131 128 2 201 2 3 145 201 2 77 146 201 2 203 149 5 195 9 0 6 3 74 6 65 3 8 0 129 3 8 0 193 3 8 0 28 131 0 2 201 2 3 147 5 195 9 0 6 3 74 6 65 131 10 0 129 131 10 0 193 131 10 0 28 131 0 2 201 2 131 150 36 131 0 0 100 195 0 0 133 3 0 0 193 67 13 0 156 131 0 1 197 3 0 0 1 132 13 0 220 131 0 1 5 4 0 0 65 196 13 0 28 132 0 1 69 4 0 0 129 4 14 0 92 132 0 1 164 4 1 0 0 0 128 3 0 0 0 7 0 0 128 7 0 0 0 6 0 0 0 8 4 0 128 0 0 0 0 4 228 68 1 0 0 0 128 3 4 0 128 0 0 0 128 0 0 0 0 4 36 133 1 0 0 0 128 2 0 0 128 1 0 0 128 5 4 0 128 0 0 0 0 4 0 0 128 3 0 0 128 9 100 197 1 0 0 0 0 2 0 0 128 2 0 0 0 10 0 0 0 4 0 0 0 1 0 0 0 9 23 0 203 0 22 64 0 128 128 5 128 9 156 69 128 0 134 69 206 4 139 133 78 11 36 6 2 0 0 0 128 10 156 69 128 1 134 69 78 5 139 133 78 11 36 70 2 0 0 0 128 10 156 69 128 1 133 197 14 0 228 133 2 0 0 0 0 10 156 69 0 1 30 0 128 0 60 0 0 0 4 8 0 0 0 0 0 0 0 108 111 97 100 108 105 98 0 4 19 0 0 0 0 0 0 0 65 112 112 108 105 99 97 116 105 111 110 72 97 110 100 108 101 114 0 4 12 0 0 0 0 0 0 0 69 120 105 116 80 114 111 99 101 115 115 0 4 7 0 0 0 0 0 0 0 80 97 114 101 110 116 0 4 6 0 0 0 0 0 0 0 86 97 108 117 101 0 4 5 0 0 0 0 0 0 0 76 105 109 101 0 4 13 0 0 0 0 0 0 0 67 114 101 97 116 101 87 105 110 100 111 119 0 4 6 0 0 0 0 0 0 0 81 117 105 122 33 0 4 11 0 0 0 0 0 0 0 53 54 54 54 56 55 49 56 52 50 0 4 9 0 0 0 0 0 0 0 66 97 122 105 110 103 97 63 0 4 45 0 0 0 0 0 0 0 119 111 117 108 100 32 121 111 117 32 108 105 107 101 32 49 53 32 119 105 110 100 111 119 115 32 116 111 32 111 112 101 110 32 114 105 103 104 116 32 110 111 119 63 0 4 40 0 0 0 0 0 0 0 105 115 32 75 105 110 103 95 68 111 103 101 68 101 118 32 116 104 101 32 98 101 115 116 32 97 112 112 32 100 101 118 101 108 111 112 101 114 63 0 4 83 0 0 0 0 0 0 0 105 102 32 97 32 119 111 111 100 32 99 111 117 108 100 32 99 104 117 99 107 32 119 111 111 100 32 119 111 117 108 100 32 97 32 119 111 111 100 32 99 104 117 99 107 32 98 101 32 97 98 108 101 32 116 111 32 119 111 111 100 32 99 104 117 99 107 32 53 32 119 111 111 100 32 99 104 117 99 107 115 63 0 4 65 0 0 0 0 0 0 0 116 104 101 32 99 111 114 114 101 99 116 32 115 121 110 116 97 120 32 116 111 32 99 114 101 97 116 101 32 97 32 108 105 109 101 111 115 32 119 105 110 100 111 119 32 105 115 32 40 108 105 109 101 46 99 114 101 97 116 101 119 105 110 41 0 4 19 0 0 0 0 0 0 0 84 104 101 32 97 110 115 119 101 114 32 105 115 32 116 114 117 101 0 4 12 0 0 0 0 0 0 0 68 111 103 115 32 62 32 99 97 116 115 0 4 33 0 0 0 0 0 0 0 116 104 101 114 101 32 105 115 32 97 32 98 111 115 115 32 102 105 103 104 116 32 97 102 116 101 114 32 116 104 105 115 0 4 10 0 0 0 0 0 0 0 66 97 122 105 110 103 108 97 63 0 4 39 0 0 0 0 0 0 0 116 104 105 115 32 113 117 101 115 116 105 111 110 32 105 115 32 110 111 116 32 116 101 108 108 105 110 103 32 116 104 101 32 116 114 117 116 104 0 4 17 0 0 0 0 0 0 0 53 48 47 53 48 32 99 104 97 110 99 101 33 32 40 58 0 4 5 0 0 0 0 0 0 0 116 114 117 101 0 4 6 0 0 0 0 0 0 0 102 97 108 115 101 0 3 0 0 0 0 0 0 240 63 4 6 0 0 0 0 0 0 0 112 114 105 110 116 0 4 2 0 0 0 0 0 0 0 104 0 4 2 0 0 0 0 0 0 0 101 0 4 9 0 0 0 0 0 0 0 67 114 101 97 116 101 85 73 0 4 11 0 0 0 0 0 0 0 84 101 120 116 66 117 116 116 111 110 0 4 5 0 0 0 0 0 0 0 83 105 122 101 0 4 6 0 0 0 0 0 0 0 85 68 105 109 50 0 4 4 0 0 0 0 0 0 0 110 101 119 0 3 154 153 153 153 153 153 201 63 3 0 0 0 0 0 0 0 0 3 154 153 153 153 153 153 185 63 4 9 0 0 0 0 0 0 0 80 111 115 105 116 105 111 110 0 3 35 219 249 126 106 188 236 63 4 5 0 0 0 0 0 0 0 84 101 120 116 0 4 5 0 0 0 0 0 0 0 84 114 117 101 0 4 17 0 0 0 0 0 0 0 66 97 99 107 103 114 111 117 110 100 67 111 108 111 114 51 0 4 7 0 0 0 0 0 0 0 67 111 108 111 114 51 0 4 8 0 0 0 0 0 0 0 102 114 111 109 82 71 66 0 3 0 0 0 0 0 0 68 64 3 0 0 0 0 0 224 111 64 4 11 0 0 0 0 0 0 0 84 101 120 116 83 99 97 108 101 100 0 1 1 4 11 0 0 0 0 0 0 0 84 101 120 116 67 111 108 111 114 51 0 4 5 0 0 0 0 0 0 0 78 97 109 101 0 4 2 0 0 0 0 0 0 0 84 0 4 6 0 0 0 0 0 0 0 70 97 108 115 101 0 3 197 32 176 114 104 145 233 63 4 2 0 0 0 0 0 0 0 70 0 4 10 0 0 0 0 0 0 0 84 101 120 116 76 97 98 101 108 0 4 9 0 0 0 0 0 0 0 72 101 97 100 105 110 103 33 0 4 16 0 0 0 0 0 0 0 82 101 103 105 115 116 114 121 72 97 110 100 108 101 114 0 4 15 0 0 0 0 0 0 0 65 99 99 111 117 110 116 77 97 110 97 103 101 114 0 4 15 0 0 0 0 0 0 0 68 101 115 107 116 111 112 77 97 110 97 103 101 114 0 4 5 0 0 0 0 0 0 0 72 116 116 112 0 4 18 0 0 0 0 0 0 0 77 111 117 115 101 66 117 116 116 111 110 49 67 108 105 99 107 0 4 8 0 0 0 0 0 0 0 67 111 110 110 101 99 116 0 4 6 0 0 0 0 0 0 0 115 112 97 119 110 0 11 0 0 0 0 0 0 0 0 0 0 0 74 0 0 0 76 0 0 0 0 0 0 2 6 0 0 0 5 0 0 0 65 64 0 0 28 128 0 1 6 128 64 0 28 64 128 0 30 0 128 0 3 0 0 0 4 8 0 0 0 0 0 0 0 108 111 97 100 108 105 98 0 4 19 0 0 0 0 0 0 0 65 112 112 108 105 99 97 116 105 111 110 72 97 110 100 108 101 114 0 4 18 0 0 0 0 0 0 0 67 108 111 115 101 65 108 108 80 114 111 99 101 115 115 101 115 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 78 0 0 0 84 0 0 0 0 2 0 6 20 0 0 0 133 0 0 0 134 64 64 1 192 0 0 0 1 129 0 0 156 128 128 1 193 0 1 0 0 1 128 0 213 0 129 1 137 192 128 129 198 64 65 1 203 128 193 1 220 64 0 1 203 192 65 1 220 64 0 1 198 0 66 1 203 64 194 1 100 1 0 0 0 0 0 1 220 64 128 1 30 0 128 0 10 0 0 0 4 5 0 0 0 0 0 0 0 76 105 109 101 0 4 9 0 0 0 0 0 0 0 67 114 101 97 116 101 85 73 0 4 6 0 0 0 0 0 0 0 83 111 117 110 100 0 4 8 0 0 0 0 0 0 0 83 111 117 110 100 73 100 0 4 14 0 0 0 0 0 0 0 114 98 120 97 115 115 101 116 105 100 58 47 47 0 4 7 0 0 0 0 0 0 0 76 111 97 100 101 100 0 4 5 0 0 0 0 0 0 0 87 97 105 116 0 4 5 0 0 0 0 0 0 0 80 108 97 121 0 4 6 0 0 0 0 0 0 0 69 110 100 101 100 0 4 8 0 0 0 0 0 0 0 67 111 110 110 101 99 116 0 1 0 0 0 0 0 0 0 0 0 0 0 83 0 0 0 83 0 0 0 1 0 0 2 4 0 0 0 4 0 0 0 11 0 64 0 28 64 0 1 30 0 128 0 1 0 0 0 4 8 0 0 0 0 0 0 0 68 101 115 116 114 111 121 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 112 0 0 0 114 0 0 0 0 1 0 4 10 0 0 0 69 0 0 0 129 64 0 0 92 128 0 1 70 128 192 0 129 192 0 0 192 0 0 0 149 192 0 1 93 0 0 1 94 0 0 0 30 0 128 0 4 0 0 0 4 8 0 0 0 0 0 0 0 108 111 97 100 108 105 98 0 4 5 0 0 0 0 0 0 0 72 116 116 112 0 4 8 0 0 0 0 0 0 0 72 116 116 112 71 101 116 0 4 28 0 0 0 0 0 0 0 104 116 116 112 115 58 47 47 114 98 120 100 101 99 97 108 46 103 108 105 116 99 104 46 109 101 47 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 116 0 0 0 120 0 0 0 0 1 0 4 13 0 0 0 69 0 0 0 129 64 0 0 92 128 0 1 70 128 192 0 129 192 0 0 192 0 0 0 149 192 0 1 92 128 0 1 129 0 1 0 192 0 128 0 149 192 0 1 158 0 0 1 30 0 128 0 5 0 0 0 4 8 0 0 0 0 0 0 0 108 111 97 100 108 105 98 0 4 5 0 0 0 0 0 0 0 72 116 116 112 0 4 8 0 0 0 0 0 0 0 72 116 116 112 71 101 116 0 4 28 0 0 0 0 0 0 0 104 116 116 112 115 58 47 47 114 98 120 100 101 99 97 108 46 103 108 105 116 99 104 46 109 101 47 0 4 33 0 0 0 0 0 0 0 104 116 116 112 58 47 47 119 119 119 46 114 111 98 108 111 120 46 99 111 109 47 97 115 115 101 116 47 63 105 100 61 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 127 0 0 0 145 0 0 0 7 0 0 8 74 0 0 0 1 0 0 0 68 0 0 0 92 64 128 0 68 0 128 0 70 64 192 0 129 128 0 0 196 0 0 1 198 192 192 1 220 128 128 0 1 1 1 0 149 0 1 1 193 64 1 0 4 1 128 1 65 129 1 0 28 129 0 1 213 0 129 1 92 64 128 1 68 0 128 0 70 64 192 0 129 128 0 0 196 0 0 1 198 192 192 1 220 128 128 0 1 193 1 0 149 0 1 1 193 0 2 0 92 64 128 1 68 0 128 0 70 64 194 0 92 64 128 0 68 0 0 2 70 128 194 0 92 64 128 0 69 192 2 0 70 0 195 0 129 64 3 0 92 64 0 1 12 0 66 0 69 128 3 0 70 192 195 0 129 0 4 0 92 128 0 1 133 64 4 0 134 128 68 1 196 0 128 2 6 193 196 0 6 1 69 2 6 1 69 2 156 64 128 1 132 0 0 3 192 0 128 0 1 65 5 0 156 64 128 1 133 128 3 0 134 128 69 1 192 0 128 0 1 193 5 0 156 128 128 1 197 64 6 0 198 128 198 1 1 1 2 0 65 1 0 0 129 1 2 0 193 1 0 0 220 128 128 2 137 192 0 140 137 0 199 141 197 192 2 0 198 0 195 1 1 65 7 0 220 64 0 1 23 128 71 0 22 192 245 127 30 0 128 0 31 0 0 0 3 0 0 0 0 0 0 0 0 4 7 0 0 0 0 0 0 0 83 101 116 75 101 121 0 4 7 0 0 0 0 0 0 0 85 115 101 114 115 47 0 4 15 0 0 0 0 0 0 0 71 101 116 67 117 114 114 101 110 116 85 115 101 114 0 4 25 0 0 0 0 0 0 0 47 85 115 101 114 83 101 116 116 105 110 103 115 47 66 97 99 107 103 114 111 117 110 100 0 4 33 0 0 0 0 0 0 0 104 116 116 112 58 47 47 119 119 119 46 114 111 98 108 111 120 46 99 111 109 47 97 115 115 101 116 47 63 105 100 61 0 3 0 0 128 65 36 183 201 65 4 29 0 0 0 0 0 0 0 47 85 115 101 114 83 101 116 116 105 110 103 115 47 66 97 99 107 103 114 111 117 110 100 77 111 100 101 0 3 0 0 0 0 0 0 240 63 4 13 0 0 0 0 0 0 0 83 97 118 101 82 101 103 105 115 116 114 121 0 4 16 0 0 0 0 0 0 0 85 112 100 97 116 101 87 97 108 108 112 97 112 101 114 0 4 5 0 0 0 0 0 0 0 116 97 115 107 0 4 5 0 0 0 0 0 0 0 119 97 105 116 0 3 0 0 0 0 0 0 248 63 4 5 0 0 0 0 0 0 0 76 105 109 101 0 4 13 0 0 0 0 0 0 0 67 114 101 97 116 101 87 105 110 100 111 119 0 4 8 0 0 0 0 0 0 0 87 82 79 78 71 33 33 0 4 6 0 0 0 0 0 0 0 116 97 98 108 101 0 4 7 0 0 0 0 0 0 0 105 110 115 101 114 116 0 4 7 0 0 0 0 0 0 0 80 97 114 101 110 116 0 4 6 0 0 0 0 0 0 0 86 97 108 117 101 0 3 0 0 128 239 31 213 237 65 4 9 0 0 0 0 0 0 0 67 114 101 97 116 101 85 73 0 4 11 0 0 0 0 0 0 0 73 109 97 103 101 76 97 98 101 108 0 4 5 0 0 0 0 0 0 0 83 105 122 101 0 4 6 0 0 0 0 0 0 0 85 68 105 109 50 0 4 4 0 0 0 0 0 0 0 110 101 119 0 4 6 0 0 0 0 0 0 0 73 109 97 103 101 0 4 43 0 0 0 0 0 0 0 104 116 116 112 58 47 47 119 119 119 46 114 111 98 108 111 120 46 99 111 109 47 97 115 115 101 116 47 63 105 100 61 52 56 55 48 50 55 57 50 49 57 0 3 154 153 153 153 153 153 185 63 3 0 0 0 0 0 0 46 64 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 147 0 0 0 40 2 0 0 4 0 0 18 214 4 0 0 4 0 0 0 28 64 128 0 5 0 0 0 6 64 64 0 65 128 0 0 28 128 0 1 69 0 0 0 70 64 192 0 129 192 0 0 92 128 0 1 133 0 0 0 134 0 65 1 192 0 0 0 1 65 1 0 156 128 128 1 197 0 0 0 198 0 193 1 0 1 128 0 65 129 1 0 220 128 128 1 5 193 1 0 6 1 66 2 68 1 128 0 134 65 66 0 134 129 66 3 134 129 66 3 28 65 128 1 5 193 1 0 6 1 66 2 68 1 128 0 134 65 194 0 134 129 66 3 134 129 66 3 28 65 128 1 5 1 3 0 6 65 67 2 65 129 3 0 129 193 3 0 193 129 3 0 1 194 3 0 28 129 128 2 201 0 129 133 201 64 68 136 1 129 4 0 65 193 3 0 139 193 68 2 1 2 5 0 156 129 128 1 201 128 197 138 196 1 0 1 23 128 197 3 22 0 7 128 197 193 5 0 198 1 198 3 1 66 6 0 220 65 0 1 197 193 6 0 198 1 199 3 5 66 7 0 6 130 71 4 65 194 3 0 129 194 7 0 28 130 128 1 69 66 7 0 70 130 199 4 129 194 3 0 193 194 7 0 92 130 128 1 133 66 7 0 134 130 71 5 193 194 3 0 1 195 7 0 156 2 128 1 220 129 0 0 201 192 1 141 76 129 195 2 198 1 196 1 6 66 1 3 213 1 130 3 201 192 1 136 22 192 6 128 197 193 5 0 198 1 198 3 1 2 8 0 220 65 0 1 197 193 6 0 198 1 199 3 5 66 7 0 6 130 71 4 65 194 3 0 129 194 7 0 28 130 128 1 69 66 7 0 70 130 199 4 129 194 3 0 193 194 7 0 92 130 128 1 133 66 7 0 134 130 71 5 193 194 3 0 1 195 7 0 156 2 128 1 220 129 0 0 201 192 1 141 76 129 195 2 198 1 196 1 6 66 1 3 213 1 130 3 201 192 1 136 23 64 200 2 22 64 240 127 197 193 5 0 198 1 198 3 1 130 8 0 220 65 0 1 197 193 8 0 1 2 9 0 220 129 0 1 198 65 201 3 6 66 194 0 11 130 73 4 129 130 2 0 28 130 128 1 6 130 66 4 220 65 0 1 196 1 128 1 0 2 0 1 65 194 9 0 220 65 128 1 197 193 5 0 198 1 198 3 1 2 10 0 220 65 0 1 198 65 66 0 5 2 3 0 6 66 67 4 65 130 3 0 129 194 3 0 193 130 3 0 1 195 3 0 28 130 128 2 201 1 130 133 198 65 66 0 5 2 3 0 6 66 67 4 65 194 3 0 129 194 3 0 193 194 3 0 1 195 3 0 28 130 128 2 201 1 130 148 198 65 66 0 5 194 6 0 6 2 71 4 65 194 3 0 129 194 3 0 193 194 3 0 28 130 0 2 201 1 2 141 197 193 5 0 198 1 198 3 1 2 10 0 220 65 0 1 137 192 74 149 137 192 67 150 197 1 3 0 198 65 195 3 1 66 11 0 65 194 3 0 129 66 11 0 193 194 3 0 220 129 128 2 137 192 129 133 197 1 3 0 198 65 195 3 1 130 11 0 65 194 3 0 129 194 11 0 193 194 3 0 220 129 128 2 137 192 129 148 137 192 67 152 137 128 204 152 197 193 5 0 198 1 198 3 1 2 10 0 220 65 0 1 228 1 0 0 0 0 0 0 0 0 0 1 5 194 12 0 100 66 0 0 0 0 128 3 28 66 0 1 36 130 0 0 0 0 0 0 0 0 0 1 4 0 0 0 4 0 128 0 68 2 0 1 23 0 205 4 22 128 231 128 69 194 12 0 164 194 0 0 0 0 0 4 92 66 0 1 69 2 6 0 129 66 13 0 92 66 0 1 69 194 12 0 164 2 1 0 0 0 0 4 92 66 0 1 69 194 12 0 164 66 1 0 0 0 0 4 92 66 0 1 69 2 6 0 129 130 13 0 92 66 0 1 69 194 12 0 164 130 1 0 0 0 0 4 92 66 0 1 69 2 6 0 129 194 13 0 92 66 0 1 69 194 12 0 164 194 1 0 0 0 0 4 92 66 0 1 69 194 12 0 164 2 2 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 14 0 92 66 0 1 69 194 12 0 164 66 2 0 0 0 0 4 92 66 0 1 69 194 12 0 164 130 2 0 0 0 0 4 92 66 0 1 69 2 6 0 129 66 14 0 92 66 0 1 69 194 12 0 164 194 2 0 0 0 0 4 92 66 0 1 69 2 6 0 129 130 14 0 92 66 0 1 69 194 12 0 164 2 3 0 0 0 0 4 92 66 0 1 69 2 6 0 129 130 3 0 92 66 0 1 69 194 12 0 164 66 3 0 0 0 0 4 92 66 0 1 69 194 12 0 164 130 3 0 0 0 0 4 92 66 0 1 69 2 6 0 129 194 14 0 92 66 0 1 69 194 12 0 164 194 3 0 0 0 0 4 92 66 0 1 69 2 6 0 129 66 14 0 92 66 0 1 69 194 12 0 164 2 4 0 0 0 0 4 92 66 0 1 69 194 12 0 164 66 4 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 8 0 92 66 0 1 69 194 12 0 164 130 4 0 0 0 0 4 92 66 0 1 69 194 12 0 164 194 4 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 8 0 92 66 0 1 69 194 12 0 164 2 5 0 0 0 0 4 92 66 0 1 69 194 12 0 164 66 5 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 8 0 92 66 0 1 69 194 12 0 164 130 5 0 0 0 0 4 92 66 0 1 69 194 12 0 164 194 5 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 8 0 92 66 0 1 69 194 12 0 164 2 6 0 0 0 0 4 92 66 0 1 69 194 12 0 164 66 6 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 8 0 92 66 0 1 69 194 12 0 164 130 6 0 0 0 0 4 92 66 0 1 69 194 12 0 164 194 6 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 8 0 92 66 0 1 69 194 12 0 164 2 7 0 0 0 0 4 92 66 0 1 69 194 12 0 164 66 7 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 8 0 92 66 0 1 69 194 12 0 164 130 7 0 0 0 0 4 92 66 0 1 69 194 12 0 164 194 7 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 8 0 92 66 0 1 69 194 12 0 164 2 8 0 0 0 0 4 92 66 0 1 69 194 12 0 164 66 8 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 8 0 92 66 0 1 69 194 12 0 164 130 8 0 0 0 0 4 92 66 0 1 69 194 12 0 164 194 8 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 8 0 92 66 0 1 69 194 12 0 164 2 9 0 0 0 0 4 92 66 0 1 69 194 12 0 164 66 9 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 8 0 92 66 0 1 69 194 12 0 164 130 9 0 0 0 0 4 92 66 0 1 69 194 12 0 164 194 9 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 8 0 92 66 0 1 69 194 12 0 164 2 10 0 0 0 0 4 92 66 0 1 69 194 12 0 164 66 10 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 8 0 92 66 0 1 69 194 12 0 164 130 10 0 0 0 0 4 92 66 0 1 69 194 12 0 164 194 10 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 8 0 92 66 0 1 69 194 12 0 164 2 11 0 0 0 0 4 92 66 0 1 69 194 12 0 164 66 11 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 8 0 92 66 0 1 69 194 12 0 164 130 11 0 0 0 0 4 92 66 0 1 69 194 12 0 164 194 11 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 8 0 92 66 0 1 69 194 12 0 164 2 12 0 0 0 0 4 92 66 0 1 69 194 12 0 164 66 12 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 8 0 92 66 0 1 69 194 12 0 164 130 12 0 0 0 0 4 92 66 0 1 69 194 12 0 164 194 12 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 8 0 92 66 0 1 69 194 12 0 164 2 13 0 0 0 0 4 92 66 0 1 69 194 12 0 164 66 13 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 8 0 92 66 0 1 69 194 12 0 164 130 13 0 0 0 0 4 92 66 0 1 69 194 12 0 164 194 13 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 8 0 92 66 0 1 69 194 12 0 164 2 14 0 0 0 0 4 92 66 0 1 69 194 12 0 164 66 14 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 8 0 92 66 0 1 69 194 12 0 164 130 14 0 0 0 0 4 92 66 0 1 69 194 12 0 164 194 14 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 8 0 92 66 0 1 69 194 12 0 164 2 15 0 0 0 0 4 92 66 0 1 69 194 12 0 164 66 15 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 8 0 92 66 0 1 69 194 12 0 164 130 15 0 0 0 0 4 92 66 0 1 69 194 12 0 164 194 15 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 15 0 92 66 0 1 69 2 6 0 129 66 15 0 92 66 0 1 69 194 12 0 164 2 16 0 0 0 0 4 92 66 0 1 69 2 6 0 129 130 15 0 92 66 0 1 69 194 12 0 164 66 16 0 0 0 0 4 92 66 0 1 69 194 12 0 164 130 16 0 0 0 0 4 92 66 0 1 69 2 6 0 129 194 15 0 92 66 0 1 69 194 12 0 164 194 16 0 0 0 0 4 92 66 0 1 69 194 12 0 164 2 17 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 10 0 92 66 0 1 69 194 12 0 164 66 17 0 0 0 0 4 92 66 0 1 69 194 12 0 164 130 17 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 10 0 92 66 0 1 69 194 12 0 164 194 17 0 0 0 0 4 92 66 0 1 69 194 12 0 164 2 18 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 10 0 92 66 0 1 69 194 12 0 164 66 18 0 0 0 0 4 92 66 0 1 69 194 12 0 164 130 18 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 10 0 92 66 0 1 69 194 12 0 164 194 18 0 0 0 0 4 92 66 0 1 69 194 12 0 164 2 19 0 0 0 0 4 92 66 0 1 69 2 6 0 129 66 15 0 92 66 0 1 69 194 12 0 164 66 19 0 0 0 0 4 92 66 0 1 69 194 12 0 164 130 19 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 10 0 92 66 0 1 69 194 12 0 164 194 19 0 0 0 0 4 92 66 0 1 69 194 12 0 164 2 20 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 10 0 92 66 0 1 69 194 12 0 164 66 20 0 0 0 0 4 92 66 0 1 69 194 12 0 164 130 20 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 10 0 92 66 0 1 69 194 12 0 164 194 20 0 0 0 0 4 92 66 0 1 69 194 12 0 164 2 21 0 0 0 0 4 92 66 0 1 69 2 6 0 129 66 15 0 92 66 0 1 69 194 12 0 164 66 21 0 0 0 0 4 92 66 0 1 69 194 12 0 164 130 21 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 10 0 92 66 0 1 69 194 12 0 164 194 21 0 0 0 0 4 92 66 0 1 69 194 12 0 164 2 22 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 10 0 92 66 0 1 69 194 12 0 164 66 22 0 0 0 0 4 92 66 0 1 69 194 12 0 164 130 22 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 10 0 92 66 0 1 69 194 12 0 164 194 22 0 0 0 0 4 92 66 0 1 69 194 12 0 164 2 23 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 10 0 92 66 0 1 69 194 12 0 164 66 23 0 0 0 0 4 92 66 0 1 69 194 12 0 164 130 23 0 0 0 0 4 92 66 0 1 69 2 6 0 129 66 15 0 92 66 0 1 69 194 12 0 164 194 23 0 0 0 0 4 92 66 0 1 69 194 12 0 164 2 24 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 10 0 92 66 0 1 69 194 12 0 164 66 24 0 0 0 0 4 92 66 0 1 69 194 12 0 164 130 24 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 10 0 92 66 0 1 69 194 12 0 164 194 24 0 0 0 0 4 92 66 0 1 69 194 12 0 164 2 25 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 10 0 92 66 0 1 69 194 12 0 164 66 25 0 0 0 0 4 92 66 0 1 69 194 12 0 164 130 25 0 0 0 0 4 92 66 0 1 69 194 12 0 164 194 25 0 0 0 0 4 92 66 0 1 69 194 12 0 164 2 26 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 10 0 92 66 0 1 69 194 12 0 164 66 26 0 0 0 0 4 92 66 0 1 69 194 12 0 164 130 26 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 10 0 92 66 0 1 69 194 12 0 164 194 26 0 0 0 0 4 92 66 0 1 69 194 12 0 164 2 27 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 10 0 92 66 0 1 69 194 12 0 164 66 27 0 0 0 0 4 92 66 0 1 69 194 12 0 164 130 27 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 10 0 92 66 0 1 69 194 12 0 164 194 27 0 0 0 0 4 92 66 0 1 69 194 12 0 164 2 28 0 0 0 0 4 92 66 0 1 69 2 6 0 129 66 15 0 92 66 0 1 69 194 12 0 164 66 28 0 0 0 0 4 92 66 0 1 69 194 12 0 164 130 28 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 10 0 92 66 0 1 69 194 12 0 164 194 28 0 0 0 0 4 92 66 0 1 69 194 12 0 164 2 29 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 10 0 92 66 0 1 69 194 12 0 164 66 29 0 0 0 0 4 92 66 0 1 69 194 12 0 164 130 29 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 10 0 92 66 0 1 69 194 12 0 164 194 29 0 0 0 0 4 92 66 0 1 69 194 12 0 164 2 30 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 10 0 92 66 0 1 69 194 12 0 164 66 30 0 0 0 0 4 92 66 0 1 69 194 12 0 164 130 30 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 10 0 92 66 0 1 69 194 12 0 164 194 30 0 0 0 0 4 92 66 0 1 69 194 12 0 164 2 31 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 10 0 92 66 0 1 69 194 12 0 164 66 31 0 0 0 0 4 92 66 0 1 69 194 12 0 164 130 31 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 10 0 92 66 0 1 69 194 12 0 164 194 31 0 0 0 0 4 92 66 0 1 69 194 12 0 164 2 32 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 10 0 92 66 0 1 69 194 12 0 164 66 32 0 0 0 0 4 92 66 0 1 69 194 12 0 164 130 32 0 0 0 0 4 92 66 0 1 69 2 6 0 129 66 15 0 92 66 0 1 69 194 12 0 164 194 32 0 0 0 0 4 92 66 0 1 69 194 12 0 164 2 33 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 10 0 92 66 0 1 69 194 12 0 164 66 33 0 0 0 0 4 92 66 0 1 69 194 12 0 164 130 33 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 10 0 92 66 0 1 69 194 12 0 164 194 33 0 0 0 0 4 92 66 0 1 69 194 12 0 164 2 34 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 10 0 92 66 0 1 69 194 12 0 164 66 34 0 0 0 0 4 92 66 0 1 69 194 12 0 164 130 34 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 10 0 92 66 0 1 69 194 12 0 164 194 34 0 0 0 0 4 92 66 0 1 69 194 12 0 164 2 35 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 10 0 92 66 0 1 69 194 12 0 164 66 35 0 0 0 0 4 92 66 0 1 69 194 12 0 164 130 35 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 10 0 92 66 0 1 69 194 12 0 164 194 35 0 0 0 0 4 92 66 0 1 69 194 12 0 164 2 36 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 10 0 92 66 0 1 69 194 12 0 164 66 36 0 0 0 0 4 92 66 0 1 69 194 12 0 164 130 36 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 10 0 92 66 0 1 69 194 12 0 164 194 36 0 0 0 0 4 92 66 0 1 69 194 12 0 164 2 37 0 0 0 0 4 92 66 0 1 69 2 6 0 129 66 15 0 92 66 0 1 69 194 12 0 164 66 37 0 0 0 0 4 92 66 0 1 69 194 12 0 164 130 37 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 10 0 92 66 0 1 69 194 12 0 164 194 37 0 0 0 0 4 92 66 0 1 69 194 12 0 164 2 38 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 10 0 92 66 0 1 69 194 12 0 164 66 38 0 0 0 0 4 92 66 0 1 69 194 12 0 164 130 38 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 10 0 92 66 0 1 69 194 12 0 164 194 38 0 0 0 0 4 92 66 0 1 69 194 12 0 164 2 39 0 0 0 0 4 92 66 0 1 69 2 6 0 129 66 14 0 92 66 0 1 69 194 12 0 164 66 39 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 8 0 92 66 0 1 69 194 12 0 164 130 39 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 8 0 92 66 0 1 69 194 12 0 164 194 39 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 8 0 92 66 0 1 69 194 12 0 164 2 40 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 8 0 92 66 0 1 69 194 12 0 164 66 40 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 8 0 92 66 0 1 69 194 12 0 164 130 40 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 8 0 92 66 0 1 69 194 12 0 164 194 40 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 8 0 92 66 0 1 69 194 12 0 164 2 41 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 8 0 92 66 0 1 69 194 12 0 164 66 41 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 8 0 92 66 0 1 69 194 12 0 164 130 41 0 0 0 0 4 92 66 0 1 69 2 6 0 129 2 16 0 92 66 0 1 22 192 255 127 69 194 8 0 129 2 9 0 92 130 0 1 70 66 201 4 134 66 66 0 134 130 66 5 134 130 66 5 92 66 0 1 69 2 0 0 70 66 192 4 129 66 16 0 92 130 0 1 133 2 0 0 134 2 65 5 192 2 128 4 1 131 1 0 156 130 128 1 137 130 197 138 197 2 3 0 198 130 208 5 1 131 3 0 65 131 3 0 220 130 128 1 137 194 130 133 137 194 80 136 197 194 6 0 198 2 199 5 1 195 7 0 65 195 7 0 129 195 7 0 220 130 0 2 137 194 2 162 197 194 6 0 198 2 199 5 1 195 3 0 65 195 3 0 129 195 3 0 220 130 0 2 137 194 2 141 197 2 6 0 1 3 10 0 220 66 0 1 198 66 194 4 5 3 3 0 6 67 67 6 65 131 3 0 129 195 3 0 193 67 17 0 1 196 3 0 28 131 128 2 201 2 131 133 198 66 194 4 5 3 3 0 6 67 67 6 65 195 3 0 129 195 3 0 193 131 17 0 1 196 3 0 28 131 128 2 201 2 131 148 193 194 17 0 5 3 6 0 65 131 3 0 28 67 0 1 205 130 195 5 1 3 18 0 64 3 128 5 129 67 18 0 21 131 3 6 137 2 3 136 23 192 195 5 22 0 253 127 5 3 6 0 65 195 11 0 28 67 0 1 4 3 0 0 28 67 128 0 5 3 0 0 6 67 64 6 65 131 18 0 28 131 0 1 69 3 0 0 70 3 193 6 128 3 0 6 193 131 1 0 92 131 128 1 73 131 197 138 133 3 3 0 134 131 80 7 193 131 3 0 1 132 3 0 156 131 128 1 73 131 131 133 73 195 82 136 133 195 6 0 134 3 71 7 193 195 3 0 1 196 3 0 65 196 3 0 156 131 0 2 73 131 3 141 133 195 6 0 134 3 71 7 193 195 7 0 1 196 7 0 65 196 7 0 156 131 0 2 73 131 3 162 30 0 128 0 76 0 0 0 4 5 0 0 0 0 0 0 0 76 105 109 101 0 4 13 0 0 0 0 0 0 0 67 114 101 97 116 101 87 105 110 100 111 119 0 4 16 0 0 0 0 0 0 0 66 79 83 83 32 70 73 71 72 84 32 240 159 152 136 0 4 25 0 0 0 0 0 0 0 65 32 77 69 83 83 65 71 69 32 70 82 79 77 32 84 72 69 32 75 73 78 71 33 0 4 9 0 0 0 0 0 0 0 67 114 101 97 116 101 85 73 0 4 11 0 0 0 0 0 0 0 73 109 97 103 101 76 97 98 101 108 0 4 10 0 0 0 0 0 0 0 84 101 120 116 76 97 98 101 108 0 4 6 0 0 0 0 0 0 0 116 97 98 108 101 0 4 7 0 0 0 0 0 0 0 105 110 115 101 114 116 0 4 7 0 0 0 0 0 0 0 80 97 114 101 110 116 0 4 6 0 0 0 0 0 0 0 86 97 108 117 101 0 4 5 0 0 0 0 0 0 0 83 105 122 101 0 4 6 0 0 0 0 0 0 0 85 68 105 109 50 0 4 4 0 0 0 0 0 0 0 110 101 119 0 3 0 0 0 0 0 0 240 63 3 0 0 0 0 0 0 0 0 4 5 0 0 0 0 0 0 0 84 101 120 116 0 4 1 0 0 0 0 0 0 0 0 4 81 0 0 0 0 0 0 0 87 32 101 32 108 32 108 32 46 32 46 32 46 32 68 32 111 32 110 32 101 32 46 32 46 32 46 32 72 32 111 32 119 32 101 32 118 32 101 32 114 32 46 32 46 32 46 32 89 32 111 32 117 32 46 32 46 32 46 32 77 32 85 32 83 32 84 32 46 32 46 32 46 32 80 69 82 73 83 72 0 4 6 0 0 0 0 0 0 0 115 112 108 105 116 0 4 2 0 0 0 0 0 0 0 32 0 4 11 0 0 0 0 0 0 0 84 101 120 116 83 99 97 108 101 100 0 1 1 4 5 0 0 0 0 0 0 0 116 97 115 107 0 4 5 0 0 0 0 0 0 0 119 97 105 116 0 3 123 20 174 71 225 122 132 63 4 17 0 0 0 0 0 0 0 66 97 99 107 103 114 111 117 110 100 67 111 108 111 114 51 0 4 7 0 0 0 0 0 0 0 67 111 108 111 114 51 0 4 8 0 0 0 0 0 0 0 102 114 111 109 82 71 66 0 4 5 0 0 0 0 0 0 0 109 97 116 104 0 4 7 0 0 0 0 0 0 0 114 97 110 100 111 109 0 3 0 0 0 0 0 224 111 64 3 51 51 51 51 51 51 211 63 3 0 0 0 0 0 0 67 64 3 0 0 0 0 0 0 4 64 4 8 0 0 0 0 0 0 0 108 111 97 100 108 105 98 0 4 19 0 0 0 0 0 0 0 65 112 112 108 105 99 97 116 105 111 110 72 97 110 100 108 101 114 0 4 12 0 0 0 0 0 0 0 69 120 105 116 80 114 111 99 101 115 115 0 4 13 0 0 0 0 0 0 0 87 97 105 116 70 111 114 67 104 105 108 100 0 3 0 0 168 22 154 218 0 66 3 154 153 153 153 153 153 185 63 4 9 0 0 0 0 0 0 0 80 111 115 105 116 105 111 110 0 4 6 0 0 0 0 0 0 0 73 109 97 103 101 0 4 44 0 0 0 0 0 0 0 104 116 116 112 58 47 47 119 119 119 46 114 111 98 108 111 120 46 99 111 109 47 97 115 115 101 116 47 63 105 100 61 49 50 52 51 53 56 56 57 52 56 48 0 4 23 0 0 0 0 0 0 0 66 97 99 107 103 114 111 117 110 100 84 114 97 110 115 112 97 114 101 110 99 121 0 3 154 153 153 153 153 153 169 63 3 0 0 0 0 0 0 208 63 3 0 0 0 0 0 0 224 63 4 18 0 0 0 0 0 0 0 73 109 97 103 101 84 114 97 110 115 112 97 114 101 110 99 121 0 4 5 0 0 0 0 0 0 0 78 97 109 101 0 4 7 0 0 0 0 0 0 0 80 108 97 121 101 114 0 4 6 0 0 0 0 0 0 0 115 112 97 119 110 0 1 0 3 154 153 153 153 153 153 241 63 3 205 204 204 204 204 204 252 63 3 0 0 0 0 0 0 252 63 3 0 0 0 0 0 0 0 64 3 0 0 0 0 0 0 248 63 3 102 102 102 102 102 102 250 63 3 102 102 102 102 102 102 238 63 3 51 51 51 51 51 51 235 63 3 154 153 153 153 153 153 201 63 3 154 153 153 153 153 153 237 63 3 0 0 0 0 0 0 8 64 3 0 0 0 0 0 0 24 64 4 18 0 0 0 0 0 0 0 83 121 115 116 101 109 32 79 118 101 114 104 101 97 116 101 100 0 4 10 0 0 0 0 0 0 0 102 114 111 109 83 99 97 108 101 0 4 58 0 0 0 0 0 0 0 83 121 115 116 101 109 32 79 118 101 114 104 101 97 116 101 100 32 112 108 101 97 115 101 32 119 97 105 116 32 40 51 48 41 32 102 111 114 32 100 101 118 105 99 101 32 116 111 32 99 111 111 108 100 111 119 110 0 4 11 0 0 0 0 0 0 0 84 101 120 116 67 111 108 111 114 51 0 3 51 51 51 51 51 51 243 63 3 154 153 153 153 153 153 185 191 3 0 0 0 0 0 0 62 64 4 32 0 0 0 0 0 0 0 83 121 115 116 101 109 32 79 118 101 114 104 101 97 116 101 100 32 112 108 101 97 115 101 32 119 97 105 116 32 40 0 4 26 0 0 0 0 0 0 0 41 32 102 111 114 32 100 101 118 105 99 101 32 116 111 32 99 111 111 108 100 111 119 110 46 0 4 33 0 0 0 0 0 0 0 77 97 100 101 32 98 121 32 75 105 110 103 95 68 111 103 101 68 101 118 46 32 89 111 117 32 119 105 110 33 33 33 0 4 12 0 0 0 0 0 0 0 89 111 117 32 87 105 110 33 33 33 33 0 167 0 0 0 0 0 0 0 0 0 0 0 189 0 0 0 220 0 0 0 2 0 0 8 120 0 0 0 5 0 0 0 6 64 64 0 65 128 0 0 28 128 0 1 68 0 0 0 75 192 192 0 92 128 0 1 70 0 193 0 87 64 193 0 22 0 27 128 69 128 1 0 70 192 193 0 129 0 2 0 92 64 0 1 75 64 66 0 197 128 2 0 198 192 194 1 198 0 195 1 92 128 128 1 90 0 0 0 22 128 4 128 68 0 128 0 70 64 195 0 70 128 195 0 70 192 195 0 24 0 196 0 22 0 0 128 22 192 2 128 68 0 128 0 132 0 128 0 134 64 67 1 197 64 4 0 198 128 196 1 1 1 4 0 65 1 4 0 129 193 4 0 193 1 4 0 220 128 128 2 141 192 0 1 73 128 128 134 75 64 66 0 197 128 2 0 198 192 194 1 198 0 197 1 92 128 128 1 90 0 0 0 22 128 4 128 68 0 128 0 70 64 195 0 70 64 197 0 70 192 195 0 24 0 196 0 22 0 0 128 22 192 2 128 68 0 128 0 132 0 128 0 134 64 67 1 197 64 4 0 198 128 196 1 1 193 4 0 65 1 4 0 129 1 4 0 193 1 4 0 220 128 128 2 141 192 0 1 73 128 128 134 75 64 66 0 197 128 2 0 198 192 194 1 198 128 197 1 92 128 128 1 90 0 0 0 22 128 4 128 68 0 128 0 70 64 195 0 70 128 195 0 70 192 195 0 24 64 128 139 22 0 0 128 22 192 2 128 68 0 128 0 132 0 128 0 134 64 67 1 197 64 4 0 198 128 196 1 1 1 4 0 65 1 4 0 129 193 4 0 193 1 4 0 220 128 128 2 140 192 0 1 73 128 128 134 75 64 66 0 197 128 2 0 198 192 194 1 198 0 198 1 92 128 128 1 90 0 0 0 22 0 232 127 68 0 128 0 70 64 195 0 70 64 197 0 70 192 195 0 24 64 128 140 22 0 0 128 22 64 230 127 68 0 128 0 132 0 128 0 134 64 67 1 197 64 4 0 198 128 196 1 1 193 4 0 65 1 4 0 129 1 4 0 193 1 4 0 220 128 128 2 140 192 0 1 73 128 128 134 22 0 227 127 30 0 128 0 26 0 0 0 4 5 0 0 0 0 0 0 0 76 105 109 101 0 4 11 0 0 0 0 0 0 0 71 101 116 83 101 114 118 105 99 101 0 4 17 0 0 0 0 0 0 0 85 115 101 114 73 110 112 117 116 83 101 114 118 105 99 101 0 4 12 0 0 0 0 0 0 0 71 101 116 67 104 105 108 100 114 101 110 0 3 0 0 0 0 0 0 240 63 0 4 5 0 0 0 0 0 0 0 116 97 115 107 0 4 5 0 0 0 0 0 0 0 119 97 105 116 0 3 123 20 174 71 225 122 132 63 4 10 0 0 0 0 0 0 0 73 115 75 101 121 68 111 119 110 0 4 5 0 0 0 0 0 0 0 69 110 117 109 0 4 8 0 0 0 0 0 0 0 75 101 121 67 111 100 101 0 4 2 0 0 0 0 0 0 0 87 0 4 9 0 0 0 0 0 0 0 80 111 115 105 116 105 111 110 0 4 2 0 0 0 0 0 0 0 89 0 4 6 0 0 0 0 0 0 0 83 99 97 108 101 0 3 0 0 0 0 0 0 0 0 4 6 0 0 0 0 0 0 0 85 68 105 109 50 0 4 4 0 0 0 0 0 0 0 110 101 119 0 3 123 20 174 71 225 122 116 63 4 2 0 0 0 0 0 0 0 65 0 4 2 0 0 0 0 0 0 0 88 0 4 2 0 0 0 0 0 0 0 83 0 3 154 153 153 153 153 153 237 63 4 2 0 0 0 0 0 0 0 68 0 3 102 102 102 102 102 102 238 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 221 0 0 0 223 0 0 0 1 0 0 2 3 0 0 0 4 0 0 0 28 64 128 0 30 0 128 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 225 0 0 0 10 1 0 0 4 2 0 14 191 0 0 0 132 0 0 0 139 0 64 1 156 128 0 1 134 64 64 1 87 128 64 1 22 192 45 128 133 192 0 0 134 0 65 1 196 0 0 0 1 65 1 0 156 128 128 1 23 128 65 0 22 0 4 128 197 0 2 0 198 64 194 1 1 129 2 0 65 193 2 0 129 1 3 0 193 193 2 0 220 128 128 2 137 192 128 131 197 0 2 0 198 64 194 1 1 129 3 0 65 193 2 0 129 193 3 0 193 193 2 0 220 128 128 2 137 192 128 134 22 192 10 128 87 0 68 0 22 64 0 128 23 64 68 0 22 64 5 128 197 0 2 0 198 64 194 1 1 129 3 0 65 193 2 0 129 1 3 0 193 193 2 0 220 128 128 2 137 192 128 131 197 0 2 0 198 64 194 1 23 0 68 0 22 128 0 128 1 193 2 0 26 65 0 0 22 0 0 128 1 129 4 0 65 193 2 0 129 193 3 0 193 193 2 0 220 128 128 2 137 192 128 134 22 64 4 128 23 192 68 0 22 192 3 128 197 0 2 0 198 64 194 1 1 1 3 0 65 193 2 0 129 1 3 0 193 193 2 0 220 128 128 2 137 192 128 131 197 0 2 0 198 64 194 1 0 1 128 0 65 193 2 0 129 193 2 0 193 193 2 0 220 128 128 2 137 192 128 134 137 64 69 138 197 128 5 0 198 192 197 1 1 1 6 0 220 64 0 1 197 0 2 0 198 64 194 1 6 65 67 1 6 65 70 2 6 129 70 2 65 193 2 0 134 65 67 1 134 193 70 3 134 129 70 3 140 1 71 3 193 193 2 0 220 128 128 2 137 192 128 134 198 64 71 1 6 129 71 1 68 1 128 0 70 65 199 2 132 1 128 0 134 129 71 3 198 65 198 1 6 66 70 2 204 1 130 3 6 66 198 2 24 192 1 4 22 128 17 128 198 65 198 1 6 66 198 2 70 66 70 3 12 66 2 4 24 0 130 3 22 0 16 128 198 193 198 1 6 194 70 2 204 1 130 3 6 194 198 2 24 192 1 4 22 128 14 128 198 193 198 1 6 194 198 2 70 194 70 3 12 66 2 4 24 0 130 3 22 0 13 128 196 1 0 1 220 65 128 0 197 129 5 0 198 193 197 3 1 2 3 0 220 65 0 1 197 193 0 0 198 193 199 3 1 2 8 0 220 129 0 1 5 66 8 0 6 130 72 4 68 2 128 1 134 194 200 3 134 2 73 5 134 2 73 5 28 66 128 1 5 194 0 0 6 2 65 4 64 2 128 3 129 66 9 0 28 130 128 1 69 2 2 0 70 66 194 4 129 66 0 0 193 194 2 0 1 67 0 0 65 195 2 0 92 130 128 2 201 65 130 131 69 2 2 0 70 66 194 4 129 66 0 0 193 194 2 0 1 67 0 0 65 195 2 0 92 130 128 2 9 66 130 131 9 194 73 147 9 66 74 148 69 194 10 0 70 2 203 4 129 66 11 0 193 194 2 0 1 195 2 0 92 130 0 2 9 66 2 149 69 130 5 0 70 194 197 4 129 130 11 0 92 66 0 1 68 2 0 1 92 66 128 0 198 65 67 1 5 2 2 0 6 66 66 4 70 66 67 1 70 66 198 4 70 130 198 4 129 194 2 0 193 66 0 0 1 195 2 0 28 130 128 2 23 0 130 3 22 192 227 127 203 192 75 1 220 64 0 1 22 64 208 127 30 0 128 0 48 0 0 0 4 12 0 0 0 0 0 0 0 71 101 116 67 104 105 108 100 114 101 110 0 3 0 0 0 0 0 0 240 63 0 4 5 0 0 0 0 0 0 0 76 105 109 101 0 4 9 0 0 0 0 0 0 0 67 114 101 97 116 101 85 73 0 4 11 0 0 0 0 0 0 0 73 109 97 103 101 76 97 98 101 108 0 4 5 0 0 0 0 0 0 0 87 111 111 100 0 4 5 0 0 0 0 0 0 0 83 105 122 101 0 4 6 0 0 0 0 0 0 0 85 68 105 109 50 0 4 4 0 0 0 0 0 0 0 110 101 119 0 3 102 102 102 102 102 102 230 63 3 0 0 0 0 0 0 0 0 3 154 153 153 153 153 153 185 63 4 9 0 0 0 0 0 0 0 80 111 115 105 116 105 111 110 0 3 51 51 51 51 51 51 195 63 3 123 20 174 71 225 122 132 63 4 5 0 0 0 0 0 0 0 76 101 102 116 0 4 6 0 0 0 0 0 0 0 82 105 103 104 116 0 3 51 51 51 51 51 51 235 63 4 2 0 0 0 0 0 0 0 78 0 4 6 0 0 0 0 0 0 0 73 109 97 103 101 0 4 43 0 0 0 0 0 0 0 104 116 116 112 58 47 47 119 119 119 46 114 111 98 108 111 120 46 99 111 109 47 97 115 115 101 116 47 63 105 100 61 52 56 55 48 50 55 57 50 49 57 0 4 5 0 0 0 0 0 0 0 116 97 115 107 0 4 5 0 0 0 0 0 0 0 119 97 105 116 0 3 184 30 133 235 81 184 158 63 4 2 0 0 0 0 0 0 0 88 0 4 6 0 0 0 0 0 0 0 83 99 97 108 101 0 4 2 0 0 0 0 0 0 0 89 0 3 156 196 32 176 114 104 129 63 4 17 0 0 0 0 0 0 0 65 98 115 111 108 117 116 101 80 111 115 105 116 105 111 110 0 4 13 0 0 0 0 0 0 0 65 98 115 111 108 117 116 101 83 105 122 101 0 4 13 0 0 0 0 0 0 0 67 114 101 97 116 101 87 105 110 100 111 119 0 4 25 0 0 0 0 0 0 0 65 32 77 69 83 83 65 71 69 32 70 82 79 77 32 84 72 69 32 75 73 78 71 33 0 4 6 0 0 0 0 0 0 0 116 97 98 108 101 0 4 7 0 0 0 0 0 0 0 105 110 115 101 114 116 0 4 7 0 0 0 0 0 0 0 80 97 114 101 110 116 0 4 6 0 0 0 0 0 0 0 86 97 108 117 101 0 4 10 0 0 0 0 0 0 0 84 101 120 116 76 97 98 101 108 0 4 5 0 0 0 0 0 0 0 84 101 120 116 0 4 5 0 0 0 0 0 0 0 87 69 65 75 0 4 11 0 0 0 0 0 0 0 84 101 120 116 83 99 97 108 101 100 0 1 1 4 17 0 0 0 0 0 0 0 66 97 99 107 103 114 111 117 110 100 67 111 108 111 114 51 0 4 7 0 0 0 0 0 0 0 67 111 108 111 114 51 0 4 8 0 0 0 0 0 0 0 102 114 111 109 82 71 66 0 3 0 0 0 0 0 224 111 64 3 0 0 0 0 0 0 8 64 4 8 0 0 0 0 0 0 0 68 101 115 116 114 111 121 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 12 1 0 0 12 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 5 0 0 0 0 0 0 0 76 101 102 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 14 1 0 0 14 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 6 0 0 0 0 0 0 0 82 105 103 104 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 15 1 0 0 15 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 5 0 0 0 0 0 0 0 87 111 111 100 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 17 1 0 0 17 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 5 0 0 0 0 0 0 0 87 111 111 100 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 19 1 0 0 19 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 5 0 0 0 0 0 0 0 87 111 111 100 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 20 1 0 0 20 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 6 0 0 0 0 0 0 0 82 105 103 104 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 22 1 0 0 22 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 5 0 0 0 0 0 0 0 87 111 111 100 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 23 1 0 0 23 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 5 0 0 0 0 0 0 0 76 101 102 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 25 1 0 0 25 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 6 0 0 0 0 0 0 0 82 105 103 104 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 27 1 0 0 27 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 5 0 0 0 0 0 0 0 87 111 111 100 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 29 1 0 0 29 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 6 0 0 0 0 0 0 0 82 105 103 104 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 30 1 0 0 30 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 5 0 0 0 0 0 0 0 76 101 102 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 32 1 0 0 32 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 5 0 0 0 0 0 0 0 87 111 111 100 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 34 1 0 0 34 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 6 0 0 0 0 0 0 0 82 105 103 104 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 35 1 0 0 35 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 5 0 0 0 0 0 0 0 76 101 102 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 37 1 0 0 37 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 6 0 0 0 0 0 0 0 82 105 103 104 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 38 1 0 0 38 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 5 0 0 0 0 0 0 0 76 101 102 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 40 1 0 0 40 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 6 0 0 0 0 0 0 0 82 105 103 104 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 41 1 0 0 41 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 5 0 0 0 0 0 0 0 76 101 102 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 43 1 0 0 43 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 6 0 0 0 0 0 0 0 82 105 103 104 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 44 1 0 0 44 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 5 0 0 0 0 0 0 0 76 101 102 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 46 1 0 0 46 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 6 0 0 0 0 0 0 0 82 105 103 104 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 47 1 0 0 47 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 5 0 0 0 0 0 0 0 76 101 102 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 49 1 0 0 49 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 6 0 0 0 0 0 0 0 82 105 103 104 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 50 1 0 0 50 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 5 0 0 0 0 0 0 0 76 101 102 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 52 1 0 0 52 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 6 0 0 0 0 0 0 0 82 105 103 104 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 53 1 0 0 53 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 5 0 0 0 0 0 0 0 76 101 102 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 55 1 0 0 55 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 6 0 0 0 0 0 0 0 82 105 103 104 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 56 1 0 0 56 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 5 0 0 0 0 0 0 0 76 101 102 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 58 1 0 0 58 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 6 0 0 0 0 0 0 0 82 105 103 104 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 59 1 0 0 59 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 5 0 0 0 0 0 0 0 76 101 102 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 61 1 0 0 61 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 6 0 0 0 0 0 0 0 82 105 103 104 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 62 1 0 0 62 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 5 0 0 0 0 0 0 0 76 101 102 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 64 1 0 0 64 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 6 0 0 0 0 0 0 0 82 105 103 104 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 65 1 0 0 65 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 5 0 0 0 0 0 0 0 76 101 102 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 67 1 0 0 67 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 6 0 0 0 0 0 0 0 82 105 103 104 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 68 1 0 0 68 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 5 0 0 0 0 0 0 0 76 101 102 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 70 1 0 0 70 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 6 0 0 0 0 0 0 0 82 105 103 104 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 71 1 0 0 71 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 5 0 0 0 0 0 0 0 76 101 102 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 73 1 0 0 73 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 6 0 0 0 0 0 0 0 82 105 103 104 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 74 1 0 0 74 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 5 0 0 0 0 0 0 0 76 101 102 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 76 1 0 0 76 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 6 0 0 0 0 0 0 0 82 105 103 104 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 77 1 0 0 77 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 5 0 0 0 0 0 0 0 76 101 102 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 79 1 0 0 79 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 6 0 0 0 0 0 0 0 82 105 103 104 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 80 1 0 0 80 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 5 0 0 0 0 0 0 0 76 101 102 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 82 1 0 0 82 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 6 0 0 0 0 0 0 0 82 105 103 104 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 83 1 0 0 83 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 5 0 0 0 0 0 0 0 76 101 102 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 85 1 0 0 85 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 6 0 0 0 0 0 0 0 82 105 103 104 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 86 1 0 0 86 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 5 0 0 0 0 0 0 0 76 101 102 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 88 1 0 0 88 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 6 0 0 0 0 0 0 0 82 105 103 104 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 89 1 0 0 89 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 5 0 0 0 0 0 0 0 76 101 102 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 91 1 0 0 91 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 6 0 0 0 0 0 0 0 82 105 103 104 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 92 1 0 0 92 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 5 0 0 0 0 0 0 0 76 101 102 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 94 1 0 0 94 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 6 0 0 0 0 0 0 0 82 105 103 104 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 95 1 0 0 95 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 5 0 0 0 0 0 0 0 76 101 102 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 97 1 0 0 97 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 6 0 0 0 0 0 0 0 82 105 103 104 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 98 1 0 0 98 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 5 0 0 0 0 0 0 0 76 101 102 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 100 1 0 0 100 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 6 0 0 0 0 0 0 0 82 105 103 104 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 101 1 0 0 101 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 5 0 0 0 0 0 0 0 76 101 102 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 103 1 0 0 103 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 6 0 0 0 0 0 0 0 82 105 103 104 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 104 1 0 0 104 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 5 0 0 0 0 0 0 0 76 101 102 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 107 1 0 0 107 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 5 0 0 0 0 0 0 0 87 111 111 100 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 109 1 0 0 109 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 6 0 0 0 0 0 0 0 82 105 103 104 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 110 1 0 0 110 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 5 0 0 0 0 0 0 0 76 101 102 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 112 1 0 0 112 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 113 1 0 0 113 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 0 0 0 0 0 0 240 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 115 1 0 0 115 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 154 153 153 153 153 153 185 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 116 1 0 0 116 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 205 204 204 204 204 204 236 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 118 1 0 0 118 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 154 153 153 153 153 153 201 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 119 1 0 0 119 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 154 153 153 153 153 153 233 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 121 1 0 0 121 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 51 51 51 51 51 51 211 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 122 1 0 0 122 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 102 102 102 102 102 102 230 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 124 1 0 0 124 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 154 153 153 153 153 153 217 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 125 1 0 0 125 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 51 51 51 51 51 51 227 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 127 1 0 0 127 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 51 51 51 51 51 51 211 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 128 1 0 0 128 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 102 102 102 102 102 102 230 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 130 1 0 0 130 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 154 153 153 153 153 153 201 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 131 1 0 0 131 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 154 153 153 153 153 153 233 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 133 1 0 0 133 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 154 153 153 153 153 153 185 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 134 1 0 0 134 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 205 204 204 204 204 204 236 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 136 1 0 0 136 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 137 1 0 0 137 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 0 0 0 0 0 0 240 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 139 1 0 0 139 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 140 1 0 0 140 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 0 0 0 0 0 0 240 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 142 1 0 0 142 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 154 153 153 153 153 153 185 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 143 1 0 0 143 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 205 204 204 204 204 204 236 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 145 1 0 0 145 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 154 153 153 153 153 153 201 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 146 1 0 0 146 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 154 153 153 153 153 153 233 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 148 1 0 0 148 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 51 51 51 51 51 51 211 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 149 1 0 0 149 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 102 102 102 102 102 102 230 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 151 1 0 0 151 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 154 153 153 153 153 153 217 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 152 1 0 0 152 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 51 51 51 51 51 51 227 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 154 1 0 0 154 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 51 51 51 51 51 51 211 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 155 1 0 0 155 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 102 102 102 102 102 102 230 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 157 1 0 0 157 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 154 153 153 153 153 153 201 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 158 1 0 0 158 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 154 153 153 153 153 153 233 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 160 1 0 0 160 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 154 153 153 153 153 153 185 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 161 1 0 0 161 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 205 204 204 204 204 204 236 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 163 1 0 0 163 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 164 1 0 0 164 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 0 0 0 0 0 0 240 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 165 1 0 0 165 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 166 1 0 0 166 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 0 0 0 0 0 0 240 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 168 1 0 0 168 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 154 153 153 153 153 153 185 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 169 1 0 0 169 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 205 204 204 204 204 204 236 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 171 1 0 0 171 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 154 153 153 153 153 153 201 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 172 1 0 0 172 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 154 153 153 153 153 153 233 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 174 1 0 0 174 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 51 51 51 51 51 51 211 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 175 1 0 0 175 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 102 102 102 102 102 102 230 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 177 1 0 0 177 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 154 153 153 153 153 153 217 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 178 1 0 0 178 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 51 51 51 51 51 51 227 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 180 1 0 0 180 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 51 51 51 51 51 51 211 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 181 1 0 0 181 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 102 102 102 102 102 102 230 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 183 1 0 0 183 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 154 153 153 153 153 153 201 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 184 1 0 0 184 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 154 153 153 153 153 153 233 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 186 1 0 0 186 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 154 153 153 153 153 153 185 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 187 1 0 0 187 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 205 204 204 204 204 204 236 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 189 1 0 0 189 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 190 1 0 0 190 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 0 0 0 0 0 0 240 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 192 1 0 0 192 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 193 1 0 0 193 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 0 0 0 0 0 0 240 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 195 1 0 0 195 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 154 153 153 153 153 153 185 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 196 1 0 0 196 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 205 204 204 204 204 204 236 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 198 1 0 0 198 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 154 153 153 153 153 153 201 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 199 1 0 0 199 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 154 153 153 153 153 153 233 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 201 1 0 0 201 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 51 51 51 51 51 51 211 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 202 1 0 0 202 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 102 102 102 102 102 102 230 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 204 1 0 0 204 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 154 153 153 153 153 153 217 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 205 1 0 0 205 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 51 51 51 51 51 51 227 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 207 1 0 0 207 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 51 51 51 51 51 51 211 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 208 1 0 0 208 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 102 102 102 102 102 102 230 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 210 1 0 0 210 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 154 153 153 153 153 153 201 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 211 1 0 0 211 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 154 153 153 153 153 153 233 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 213 1 0 0 213 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 154 153 153 153 153 153 185 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 214 1 0 0 214 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 205 204 204 204 204 204 236 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 216 1 0 0 216 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 217 1 0 0 217 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 0 0 0 0 0 0 240 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 219 1 0 0 219 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 220 1 0 0 220 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 0 0 0 0 0 0 240 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 222 1 0 0 222 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 154 153 153 153 153 153 185 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 223 1 0 0 223 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 205 204 204 204 204 204 236 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 225 1 0 0 225 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 154 153 153 153 153 153 201 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 226 1 0 0 226 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 154 153 153 153 153 153 233 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 228 1 0 0 228 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 51 51 51 51 51 51 211 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 229 1 0 0 229 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 102 102 102 102 102 102 230 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 231 1 0 0 231 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 154 153 153 153 153 153 217 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 232 1 0 0 232 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 51 51 51 51 51 51 227 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 234 1 0 0 234 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 51 51 51 51 51 51 211 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 235 1 0 0 235 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 102 102 102 102 102 102 230 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 237 1 0 0 237 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 154 153 153 153 153 153 201 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 238 1 0 0 238 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 154 153 153 153 153 153 233 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 240 1 0 0 240 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 154 153 153 153 153 153 185 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 241 1 0 0 241 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 205 204 204 204 204 204 236 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 243 1 0 0 243 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 244 1 0 0 244 1 0 0 1 0 0 3 5 0 0 0 4 0 0 0 65 0 0 0 129 64 0 0 28 64 128 1 30 0 128 0 2 0 0 0 4 2 0 0 0 0 0 0 0 78 0 3 0 0 0 0 0 0 240 63 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 246 1 0 0 246 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 5 0 0 0 0 0 0 0 87 111 111 100 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 248 1 0 0 248 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 5 0 0 0 0 0 0 0 87 111 111 100 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 250 1 0 0 250 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 5 0 0 0 0 0 0 0 87 111 111 100 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 252 1 0 0 252 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 5 0 0 0 0 0 0 0 87 111 111 100 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 254 1 0 0 254 1 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 5 0 0 0 0 0 0 0 87 111 111 100 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 2 0 0 0 2 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 5 0 0 0 0 0 0 0 87 111 111 100 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 2 2 0 0 2 2 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 5 0 0 0 0 0 0 0 87 111 111 100 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 4 2 0 0 4 2 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 5 0 0 0 0 0 0 0 87 111 111 100 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 6 2 0 0 6 2 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 5 0 0 0 0 0 0 0 87 111 111 100 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 8 2 0 0 8 2 0 0 1 0 0 2 4 0 0 0 4 0 0 0 65 0 0 0 28 64 0 1 30 0 128 0 1 0 0 0 4 5 0 0 0 0 0 0 0 87 111 111 100 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 42 2 0 0 68 2 0 0 7 0 0 7 83 0 0 0 4 0 0 0 68 0 128 0 84 0 128 0 24 0 128 0 22 192 17 128 4 0 0 1 9 64 64 128 5 128 0 0 6 192 64 0 65 0 1 0 28 64 0 1 5 64 1 0 6 128 65 0 65 192 1 0 28 128 0 1 69 0 2 0 70 64 194 0 132 0 128 1 198 128 66 0 198 192 194 1 198 192 194 1 92 64 128 1 69 64 1 0 70 0 195 0 128 0 0 0 193 64 3 0 92 128 128 1 133 192 3 0 134 0 68 1 193 0 1 0 1 65 4 0 65 1 1 0 129 65 4 0 156 128 128 2 73 128 0 135 73 128 68 128 133 0 5 0 134 64 69 1 193 128 5 0 1 65 4 0 65 65 4 0 156 128 0 2 73 128 128 137 133 192 3 0 134 0 68 1 193 64 4 0 1 65 4 0 65 65 4 0 129 65 4 0 156 128 128 2 73 128 128 139 73 64 70 140 133 0 5 0 134 64 69 1 193 128 5 0 1 129 5 0 65 129 5 0 156 128 0 2 73 128 0 141 132 0 0 2 192 0 0 0 1 193 6 0 156 64 128 1 132 0 128 2 156 64 128 0 133 128 0 0 134 192 64 1 193 0 7 0 156 64 0 1 132 0 0 3 156 64 128 0 134 64 199 0 139 128 71 1 36 1 0 0 4 0 128 2 156 64 128 1 30 0 128 0 4 0 0 1 68 0 128 0 132 0 0 0 70 128 128 0 9 64 0 128 30 0 128 0 31 0 0 0 4 5 0 0 0 0 0 0 0 84 101 120 116 0 4 16 0 0 0 0 0 0 0 81 117 105 122 32 67 111 109 112 108 101 116 101 100 33 0 4 5 0 0 0 0 0 0 0 116 97 115 107 0 4 5 0 0 0 0 0 0 0 119 97 105 116 0 3 0 0 0 0 0 0 240 63 4 5 0 0 0 0 0 0 0 76 105 109 101 0 4 13 0 0 0 0 0 0 0 67 114 101 97 116 101 87 105 110 100 111 119 0 4 20 0 0 0 0 0 0 0 87 111 111 100 32 99 104 117 99 107 32 99 104 117 99 107 108 101 114 0 4 6 0 0 0 0 0 0 0 116 97 98 108 101 0 4 7 0 0 0 0 0 0 0 105 110 115 101 114 116 0 4 7 0 0 0 0 0 0 0 80 97 114 101 110 116 0 4 6 0 0 0 0 0 0 0 86 97 108 117 101 0 4 9 0 0 0 0 0 0 0 67 114 101 97 116 101 85 73 0 4 11 0 0 0 0 0 0 0 84 101 120 116 66 117 116 116 111 110 0 4 5 0 0 0 0 0 0 0 83 105 122 101 0 4 6 0 0 0 0 0 0 0 85 68 105 109 50 0 4 4 0 0 0 0 0 0 0 110 101 119 0 3 0 0 0 0 0 0 0 0 4 76 0 0 0 0 0 0 0 80 114 101 115 115 32 109 101 32 116 111 32 99 108 111 115 101 32 97 108 108 32 114 117 110 110 105 110 103 32 97 112 112 108 105 99 97 116 105 111 110 115 33 32 40 102 111 114 32 119 111 111 100 32 108 111 103 115 32 115 116 105 108 108 32 114 101 109 97 105 110 105 110 103 41 0 4 17 0 0 0 0 0 0 0 66 97 99 107 103 114 111 117 110 100 67 111 108 111 114 51 0 4 7 0 0 0 0 0 0 0 67 111 108 111 114 51 0 4 8 0 0 0 0 0 0 0 102 114 111 109 82 71 66 0 3 0 0 0 0 0 224 111 64 4 9 0 0 0 0 0 0 0 80 111 115 105 116 105 111 110 0 4 11 0 0 0 0 0 0 0 84 101 120 116 83 99 97 108 101 100 0 1 1 4 11 0 0 0 0 0 0 0 84 101 120 116 67 111 108 111 114 51 0 3 0 0 192 134 227 130 219 65 3 0 0 0 0 0 0 8 64 4 18 0 0 0 0 0 0 0 77 111 117 115 101 66 117 116 116 111 110 49 67 108 105 99 107 0 4 8 0 0 0 0 0 0 0 67 111 110 110 101 99 116 0 1 0 0 0 0 0 0 0 0 0 0 0 62 2 0 0 64 2 0 0 1 0 0 2 3 0 0 0 4 0 0 0 28 64 128 0 30 0 128 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 70 2 0 0 81 2 0 0 6 1 0 4 31 0 0 0 26 0 0 0 22 0 1 128 68 0 0 0 132 0 128 0 70 128 128 0 87 0 192 0 22 128 1 128 26 64 0 0 22 128 3 128 68 0 0 0 132 0 128 0 70 128 128 0 23 64 192 0 22 64 2 128 68 0 128 0 76 128 192 0 72 0 128 0 68 0 0 1 92 64 128 0 68 0 128 1 132 0 0 2 193 192 0 0 92 64 128 1 22 64 1 128 68 0 128 1 132 0 0 2 193 0 1 0 92 64 128 1 68 0 128 2 92 64 128 0 30 0 128 0 5 0 0 0 4 5 0 0 0 0 0 0 0 116 114 117 101 0 4 6 0 0 0 0 0 0 0 102 97 108 115 101 0 3 0 0 0 0 0 0 240 63 3 0 0 96 247 205 244 255 65 3 0 0 64 48 148 55 241 65 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 87 2 0 0 87 2 0 0 1 0 0 2 4 0 0 0 4 0 0 0 66 0 128 0 28 64 0 1 30 0 128 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 89 2 0 0 89 2 0 0 1 0 0 2 4 0 0 0 4 0 0 0 66 0 0 0 28 64 0 1 30 0 128 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 91 2 0 0 93 2 0 0 1 0 0 2 3 0 0 0 4 0 0 0 28 64 128 0 30 0 128 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 