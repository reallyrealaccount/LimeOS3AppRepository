76 69 70 0 0 0 0 0 1 0 0 0 0 0 0 0 57 66 105 116 66 121 116 101 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 56 57 49 101 51 54 54 97 101 99 50 99 55 48 100 52 48 53 55 51 100 50 52 55 102 53 48 100 98 49 100 98 50 55 102 98 54 99 51 48 50 98 49 102 48 54 99 102 51 56 53 54 102 98 56 48 97 98 54 49 102 51 51 101 27 76 117 97 81 0 1 4 8 4 8 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 2 56 203 2 0 0 5 0 0 0 6 64 64 0 65 128 0 0 28 128 0 1 67 0 128 0 133 0 0 0 134 192 64 1 193 0 1 0 0 1 0 0 156 128 128 1 197 128 1 0 198 192 193 1 1 1 2 0 65 1 2 0 220 128 128 1 137 192 128 130 197 128 1 0 198 192 193 1 1 129 2 0 65 129 2 0 220 128 128 1 137 192 128 132 137 0 195 133 137 128 195 134 137 0 196 135 197 128 4 0 198 192 196 1 1 1 5 0 65 1 5 0 129 1 5 0 220 128 0 2 137 192 128 136 137 128 197 138 197 0 0 0 198 192 192 1 1 193 5 0 64 1 0 0 220 128 128 1 5 129 1 0 6 193 65 2 65 1 4 0 129 1 4 0 28 129 128 1 201 0 129 130 201 64 70 140 5 1 0 0 6 193 64 2 65 193 5 0 128 1 128 1 28 129 128 1 69 129 1 0 70 193 193 2 129 129 2 0 193 129 2 0 92 129 128 1 9 65 129 130 69 129 1 0 70 193 193 2 129 129 6 0 193 129 6 0 92 129 128 1 9 65 129 132 69 129 4 0 70 193 196 2 129 1 5 0 193 1 5 0 1 2 5 0 92 129 0 2 9 65 129 141 9 65 71 142 9 65 70 140 9 129 199 138 69 1 0 0 70 193 192 2 129 1 1 0 192 1 0 2 92 129 128 1 133 129 1 0 134 193 65 3 193 65 7 0 1 194 7 0 156 129 128 1 73 129 129 130 133 129 1 0 134 193 65 3 193 1 8 0 1 2 5 0 156 129 128 1 73 129 129 132 73 1 195 133 73 65 200 134 73 1 196 135 133 129 4 0 134 193 68 3 193 129 8 0 1 130 8 0 65 130 8 0 156 129 0 2 73 129 129 136 133 1 0 0 134 193 64 3 193 193 8 0 0 2 0 2 156 129 128 1 197 129 1 0 198 193 193 3 1 2 9 0 65 2 8 0 220 129 128 1 137 193 129 130 197 129 1 0 198 193 193 3 1 194 7 0 65 194 7 0 220 129 128 1 137 193 129 132 137 1 195 133 137 65 201 134 137 129 201 135 197 129 4 0 198 193 196 3 1 130 8 0 65 130 8 0 129 130 8 0 220 129 0 2 137 193 129 136 197 1 0 0 198 193 192 3 1 194 8 0 64 2 0 2 220 129 128 1 5 130 1 0 6 194 65 4 65 2 9 0 129 2 8 0 28 130 128 1 201 1 130 130 5 130 1 0 6 194 65 4 65 194 7 0 129 194 9 0 28 130 128 1 201 1 130 132 201 1 195 133 201 1 202 134 201 129 201 135 5 130 4 0 6 194 68 4 65 130 8 0 129 130 8 0 193 130 8 0 28 130 0 2 201 1 130 136 5 2 0 0 6 194 64 4 65 194 8 0 128 2 0 2 28 130 128 1 69 130 1 0 70 194 193 4 129 2 9 0 193 2 8 0 92 130 128 1 9 66 130 130 69 130 1 0 70 194 193 4 129 194 7 0 193 66 10 0 92 130 128 1 9 66 130 132 9 2 195 133 9 130 202 134 9 130 201 135 69 130 4 0 70 194 196 4 129 130 8 0 193 130 8 0 1 131 8 0 92 130 0 2 9 66 130 136 69 2 0 0 70 194 192 4 129 194 5 0 192 2 0 0 92 130 128 1 133 130 1 0 134 194 65 5 193 2 4 0 1 3 4 0 156 130 128 1 73 130 130 130 133 2 0 0 134 194 64 5 193 194 5 0 0 3 0 0 156 130 128 1 197 130 1 0 198 194 193 5 1 3 4 0 65 3 4 0 220 130 128 1 137 194 130 130 137 66 70 140 197 2 0 0 198 194 192 5 1 195 10 0 64 3 0 5 220 130 128 1 201 2 203 134 201 130 203 150 5 131 1 0 6 195 65 6 65 67 7 0 129 3 8 0 28 131 128 1 201 2 131 130 5 131 1 0 6 195 65 6 65 3 8 0 129 131 6 0 28 131 128 1 201 2 131 132 5 3 0 0 6 195 64 6 65 195 5 0 128 3 0 0 28 131 128 1 69 131 1 0 70 195 193 6 129 3 4 0 193 3 4 0 92 131 128 1 9 67 131 130 9 67 70 140 69 3 0 0 70 195 192 6 129 195 5 0 192 3 0 0 92 131 128 1 133 131 1 0 134 195 65 7 193 3 4 0 1 4 4 0 156 131 128 1 73 131 131 130 73 67 70 140 133 3 0 0 134 195 64 7 193 3 1 0 0 4 128 6 156 131 128 1 197 131 1 0 198 195 193 7 1 68 7 0 65 196 7 0 220 131 128 1 137 195 131 130 197 131 1 0 198 195 193 7 1 4 8 0 65 4 5 0 220 131 128 1 137 195 131 132 137 3 195 133 137 195 203 134 137 3 196 135 197 131 4 0 198 195 196 7 1 132 8 0 65 132 8 0 129 132 8 0 220 131 0 2 137 195 131 136 197 3 0 0 198 195 192 7 1 196 10 0 64 4 0 6 220 131 128 1 5 132 1 0 6 196 65 8 65 68 7 0 129 196 7 0 28 132 128 1 201 3 132 130 5 132 1 0 6 196 65 8 65 4 8 0 129 4 5 0 28 132 128 1 201 3 132 132 201 3 195 133 201 3 204 134 201 67 199 135 5 132 4 0 6 196 68 8 65 132 8 0 129 132 8 0 193 132 8 0 28 132 0 2 201 3 132 136 5 4 0 0 6 196 64 8 65 196 8 0 128 4 0 5 28 132 128 1 69 132 1 0 70 196 193 8 129 4 9 0 193 4 8 0 92 132 128 1 9 68 132 130 69 132 1 0 70 196 193 8 129 196 7 0 193 68 10 0 92 132 128 1 9 68 132 132 9 4 195 133 9 68 204 134 9 132 201 135 69 132 4 0 70 196 196 8 129 132 8 0 193 132 8 0 1 133 8 0 92 132 0 2 9 68 132 136 69 4 0 0 70 196 192 8 129 132 12 0 192 4 128 4 92 132 128 1 133 132 1 0 134 196 65 9 193 4 4 0 1 5 4 0 156 132 128 1 73 132 132 130 73 4 196 135 73 4 205 153 133 4 0 0 134 196 64 9 193 4 1 0 0 5 128 4 156 132 128 1 197 132 1 0 198 196 193 9 1 69 7 0 65 197 7 0 220 132 128 1 137 196 132 130 197 132 1 0 198 196 193 9 1 5 8 0 65 5 5 0 220 132 128 1 137 196 132 132 137 4 195 133 137 132 192 134 137 4 196 135 197 132 4 0 198 196 196 9 1 133 8 0 65 133 8 0 129 133 8 0 220 132 0 2 137 196 132 136 197 4 0 0 198 196 192 9 1 197 8 0 64 5 128 4 220 132 128 1 5 133 1 0 6 197 65 10 65 5 9 0 129 5 8 0 28 133 128 1 201 4 133 130 5 133 1 0 6 197 65 10 65 197 7 0 129 197 7 0 28 133 128 1 201 4 133 132 201 4 195 133 201 68 205 134 201 132 201 135 5 133 4 0 6 197 68 10 65 133 8 0 129 133 8 0 193 133 8 0 28 133 0 2 201 4 133 136 5 5 0 0 6 197 64 10 65 197 8 0 128 5 128 4 28 133 128 1 69 133 1 0 70 197 193 10 129 5 9 0 193 5 8 0 92 133 128 1 9 69 133 130 69 133 1 0 70 197 193 10 129 197 7 0 193 197 9 0 92 133 128 1 9 69 133 132 9 5 195 133 9 5 202 134 9 133 201 135 69 133 4 0 70 197 196 10 129 133 8 0 193 133 8 0 1 134 8 0 92 133 0 2 9 69 133 136 69 5 0 0 70 197 192 10 129 197 8 0 192 5 128 4 92 133 128 1 133 133 1 0 134 197 65 11 193 5 9 0 1 6 8 0 156 133 128 1 73 133 133 130 133 133 1 0 134 197 65 11 193 197 7 0 1 70 10 0 156 133 128 1 73 133 133 132 73 5 195 133 73 133 205 134 73 133 201 135 133 133 4 0 134 197 68 11 193 133 8 0 1 134 8 0 65 134 8 0 156 133 0 2 73 133 133 136 134 197 205 10 139 5 78 11 36 6 0 0 0 0 0 0 156 69 128 1 134 197 77 10 139 5 78 11 36 70 0 0 0 0 128 4 0 0 128 1 0 0 128 6 0 0 0 5 156 69 128 1 134 197 77 8 139 5 78 11 36 134 0 0 0 0 128 6 0 0 0 5 0 0 0 2 0 0 128 4 0 0 128 1 156 69 128 1 134 197 205 3 139 5 78 11 36 198 0 0 0 0 128 4 0 0 128 1 0 0 128 6 0 0 0 5 156 69 128 1 133 5 0 0 134 197 64 11 193 69 14 0 0 6 128 1 156 133 128 1 197 133 1 0 198 197 193 11 1 6 4 0 65 6 4 0 220 133 128 1 137 197 133 130 197 133 4 0 198 197 196 11 1 6 11 0 65 6 11 0 129 6 11 0 220 133 0 2 137 197 5 157 198 197 206 5 203 5 206 11 100 6 1 0 0 0 0 11 0 0 128 5 220 69 128 1 197 5 0 0 198 197 192 11 1 6 15 0 64 6 0 11 220 133 128 1 5 6 0 0 6 198 64 12 65 70 15 0 128 6 128 11 28 134 128 1 69 6 0 0 70 198 192 12 129 6 1 0 192 6 128 1 92 134 128 1 133 134 1 0 134 198 65 13 193 6 2 0 1 7 2 0 156 134 128 1 73 134 134 130 73 134 207 134 73 6 195 133 133 134 4 0 134 198 68 13 193 134 8 0 1 135 8 0 65 135 8 0 156 134 0 2 73 134 134 136 73 6 196 135 133 134 1 0 134 198 65 13 193 198 15 0 1 199 15 0 156 134 128 1 73 134 134 132 133 6 0 0 134 198 64 13 193 6 1 0 0 7 128 1 156 134 128 1 197 134 1 0 198 198 193 13 1 7 2 0 65 7 2 0 220 134 128 1 137 198 134 130 137 6 195 133 137 6 196 135 197 134 4 0 198 198 196 13 1 7 5 0 65 7 5 0 129 7 5 0 220 134 0 2 137 198 134 136 137 6 208 134 193 6 11 0 1 7 11 0 65 71 16 0 129 135 16 0 193 199 16 0 36 72 1 0 0 0 128 14 0 0 0 12 100 136 1 0 0 0 128 14 0 0 0 15 0 0 128 15 0 0 0 16 129 200 16 0 228 200 1 0 0 0 0 14 0 0 128 13 0 0 0 17 0 0 128 16 0 0 0 7 5 9 0 0 6 201 64 18 65 9 17 0 128 9 128 11 28 137 128 1 137 5 137 162 9 201 81 163 65 9 5 0 129 9 5 0 193 9 18 0 5 10 0 0 6 74 82 20 65 138 18 0 28 138 0 1 69 202 18 0 92 138 128 0 164 10 2 0 0 0 0 20 0 0 128 18 0 0 128 19 0 0 0 19 0 0 0 18 135 10 19 0 142 74 135 166 197 10 0 0 198 202 192 21 1 203 8 0 64 11 128 1 220 138 128 1 201 138 211 138 201 10 196 135 201 202 211 134 5 139 1 0 6 203 65 22 65 11 4 0 129 11 4 0 28 139 128 1 201 10 139 130 6 203 205 21 11 11 78 22 164 75 2 0 0 0 0 20 0 0 128 11 0 0 0 18 0 0 0 21 28 75 128 1 6 11 212 21 11 11 78 22 164 139 2 0 0 0 128 11 0 0 0 18 0 0 0 21 0 0 128 14 0 0 0 16 28 75 128 1 1 75 20 0 67 11 128 22 134 139 84 20 139 11 78 23 36 204 2 0 0 0 128 1 0 0 0 20 0 0 0 2 0 0 128 21 156 139 128 1 64 11 0 23 134 203 77 3 139 11 78 23 36 12 3 0 0 0 0 20 0 0 128 21 0 0 0 2 156 75 128 1 134 203 77 4 139 11 78 23 36 76 3 0 0 0 0 12 0 0 128 11 0 0 128 0 0 0 128 1 0 0 0 2 0 0 128 4 156 75 128 1 134 203 212 20 139 11 78 23 5 12 19 0 156 75 128 1 129 11 21 0 228 139 3 0 0 0 0 18 0 0 128 14 0 0 0 23 0 0 128 11 1 12 5 0 65 76 21 0 130 12 0 0 193 140 21 0 36 205 3 0 0 0 128 0 0 0 0 20 0 0 0 18 0 0 128 23 0 0 0 22 0 0 128 11 0 0 128 14 0 0 0 23 0 0 0 24 0 0 0 25 0 0 128 24 0 0 128 25 0 0 0 13 70 205 205 9 75 13 206 26 228 13 4 0 0 0 128 4 0 0 128 1 0 0 128 6 0 0 0 5 0 0 128 17 0 0 0 18 0 0 0 20 0 0 0 26 92 77 128 1 69 205 21 0 129 13 22 0 92 141 0 1 70 77 214 26 134 141 86 0 134 205 86 27 134 205 86 27 228 77 4 0 0 0 128 0 0 0 128 22 92 77 128 1 30 0 128 0 92 0 0 0 4 5 0 0 0 0 0 0 0 76 105 109 101 0 4 13 0 0 0 0 0 0 0 67 114 101 97 116 101 87 105 110 100 111 119 0 4 11 0 0 0 0 0 0 0 66 117 105 108 100 66 114 101 97 107 0 4 9 0 0 0 0 0 0 0 67 114 101 97 116 101 85 73 0 4 10 0 0 0 0 0 0 0 84 101 120 116 76 97 98 101 108 0 4 5 0 0 0 0 0 0 0 83 105 122 101 0 4 6 0 0 0 0 0 0 0 85 68 105 109 50 0 4 10 0 0 0 0 0 0 0 102 114 111 109 83 99 97 108 101 0 3 154 153 153 153 153 153 185 63 4 9 0 0 0 0 0 0 0 80 111 115 105 116 105 111 110 0 3 205 204 204 204 204 204 236 63 4 11 0 0 0 0 0 0 0 84 101 120 116 83 99 97 108 101 100 0 1 1 4 5 0 0 0 0 0 0 0 84 101 120 116 0 4 11 0 0 0 0 0 0 0 118 48 46 49 46 48 32 100 101 118 0 4 23 0 0 0 0 0 0 0 66 97 99 107 103 114 111 117 110 100 84 114 97 110 115 112 97 114 101 110 99 121 0 3 0 0 0 0 0 0 240 63 4 11 0 0 0 0 0 0 0 84 101 120 116 67 111 108 111 114 51 0 4 7 0 0 0 0 0 0 0 67 111 108 111 114 51 0 4 8 0 0 0 0 0 0 0 102 114 111 109 82 71 66 0 3 0 0 0 0 0 0 0 0 4 7 0 0 0 0 0 0 0 90 73 110 100 101 120 0 3 0 0 0 0 0 0 38 64 4 6 0 0 0 0 0 0 0 70 114 97 109 101 0 4 8 0 0 0 0 0 0 0 86 105 115 105 98 108 101 0 1 0 3 154 153 153 153 153 153 169 63 4 17 0 0 0 0 0 0 0 66 97 99 107 103 114 111 117 110 100 67 111 108 111 114 51 0 4 13 0 0 0 0 0 0 0 84 114 97 110 115 112 97 114 101 110 99 121 0 3 51 51 51 51 51 51 227 63 3 0 0 0 0 0 0 36 64 3 51 51 51 51 51 51 211 63 3 154 153 153 153 153 153 201 63 4 7 0 0 0 0 0 0 0 80 97 117 115 101 100 0 3 0 0 0 0 0 224 111 64 4 11 0 0 0 0 0 0 0 84 101 120 116 66 117 116 116 111 110 0 3 154 153 153 153 153 153 217 63 4 13 0 0 0 0 0 0 0 66 97 99 107 32 116 111 32 103 97 109 101 0 3 102 102 102 102 102 102 230 63 3 205 204 204 204 204 204 224 63 4 9 0 0 0 0 0 0 0 83 101 116 116 105 110 103 115 0 3 0 0 0 0 0 0 232 63 4 15 0 0 0 0 0 0 0 82 101 116 117 114 110 32 116 111 32 109 101 110 117 0 4 8 0 0 0 0 0 0 0 84 101 120 116 66 111 120 0 3 0 0 0 0 0 0 89 64 4 16 0 0 0 0 0 0 0 80 108 97 99 101 104 111 108 100 101 114 84 101 120 116 0 4 6 0 0 0 0 0 0 0 48 45 50 53 53 0 4 11 0 0 0 0 0 0 0 76 111 97 100 105 110 103 46 46 46 0 4 5 0 0 0 0 0 0 0 83 101 101 100 0 4 5 0 0 0 0 0 0 0 66 97 99 107 0 4 11 0 0 0 0 0 0 0 73 109 97 103 101 76 97 98 101 108 0 4 6 0 0 0 0 0 0 0 73 109 97 103 101 0 4 43 0 0 0 0 0 0 0 104 116 116 112 58 47 47 119 119 119 46 114 111 98 108 111 120 46 99 111 109 47 97 115 115 101 116 47 63 105 100 61 56 50 55 53 50 48 57 54 54 48 0 4 6 0 0 0 0 0 0 0 80 108 97 121 33 0 4 5 0 0 0 0 0 0 0 81 117 105 116 0 4 18 0 0 0 0 0 0 0 77 111 117 115 101 66 117 116 116 111 110 49 67 108 105 99 107 0 4 8 0 0 0 0 0 0 0 67 111 110 110 101 99 116 0 4 14 0 0 0 0 0 0 0 86 105 101 119 112 111 114 116 70 114 97 109 101 0 4 8 0 0 0 0 0 0 0 65 109 98 105 101 110 116 0 4 10 0 0 0 0 0 0 0 70 111 99 117 115 76 111 115 116 0 4 11 0 0 0 0 0 0 0 87 111 114 108 100 77 111 100 101 108 0 4 7 0 0 0 0 0 0 0 70 111 108 100 101 114 0 4 2 0 0 0 0 0 0 0 43 0 3 205 204 204 204 204 204 220 63 4 4 0 0 0 0 0 0 0 70 80 83 0 3 0 0 0 0 0 0 0 64 3 0 0 0 0 0 0 78 64 3 0 0 0 0 0 0 68 64 4 7 0 0 0 0 0 0 0 67 97 109 101 114 97 0 4 14 0 0 0 0 0 0 0 67 117 114 114 101 110 116 67 97 109 101 114 97 0 4 11 0 0 0 0 0 0 0 67 97 109 101 114 97 84 121 112 101 0 4 11 0 0 0 0 0 0 0 83 99 114 105 112 116 97 98 108 101 0 3 0 0 0 0 0 0 224 191 4 11 0 0 0 0 0 0 0 71 101 116 83 101 114 118 105 99 101 0 4 17 0 0 0 0 0 0 0 85 115 101 114 73 110 112 117 116 83 101 114 118 105 99 101 0 4 9 0 0 0 0 0 0 0 71 101 116 77 111 117 115 101 0 4 10 0 0 0 0 0 0 0 77 111 117 115 101 77 111 118 101 0 3 0 0 0 0 0 0 20 64 3 0 0 0 0 0 56 143 64 4 1 0 0 0 0 0 0 0 0 4 18 0 0 0 0 0 0 0 77 111 117 115 101 66 117 116 116 111 110 50 67 108 105 99 107 0 3 0 0 0 0 0 0 224 63 4 11 0 0 0 0 0 0 0 73 110 112 117 116 66 101 103 97 110 0 4 5 0 0 0 0 0 0 0 77 111 118 101 0 3 123 20 174 71 225 122 132 63 3 120 170 221 16 68 119 226 191 3 154 153 153 153 153 153 233 63 4 8 0 0 0 0 0 0 0 108 111 97 100 108 105 98 0 4 19 0 0 0 0 0 0 0 65 112 112 108 105 99 97 116 105 111 110 72 97 110 100 108 101 114 0 4 7 0 0 0 0 0 0 0 79 110 69 120 105 116 0 4 7 0 0 0 0 0 0 0 80 97 114 101 110 116 0 4 6 0 0 0 0 0 0 0 86 97 108 117 101 0 18 0 0 0 0 0 0 0 0 0 0 0 140 0 0 0 142 0 0 0 1 0 0 2 9 0 0 0 5 0 0 0 65 64 0 0 28 128 0 1 6 128 64 0 6 192 64 0 68 0 0 0 70 0 193 0 28 64 0 1 30 0 128 0 5 0 0 0 4 8 0 0 0 0 0 0 0 108 111 97 100 108 105 98 0 4 19 0 0 0 0 0 0 0 65 112 112 108 105 99 97 116 105 111 110 72 97 110 100 108 101 114 0 4 5 0 0 0 0 0 0 0 85 115 101 114 0 4 10 0 0 0 0 0 0 0 67 108 111 115 101 80 114 111 99 0 4 7 0 0 0 0 0 0 0 80 97 114 101 110 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 144 0 0 0 149 0 0 0 4 0 0 2 9 0 0 0 4 0 0 0 9 64 64 128 4 0 128 0 9 64 64 128 4 0 0 1 9 64 64 128 4 0 128 1 9 128 64 128 30 0 128 0 3 0 0 0 4 8 0 0 0 0 0 0 0 86 105 115 105 98 108 101 0 1 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 151 0 0 0 161 0 0 0 5 0 0 2 18 0 0 0 4 0 0 0 9 64 64 128 4 0 128 0 9 64 64 128 4 0 0 1 6 0 64 0 26 0 0 0 22 0 1 128 4 0 128 1 9 64 64 128 4 0 0 2 9 128 64 128 22 192 0 128 4 0 128 1 9 128 64 128 4 0 0 2 9 64 64 128 30 0 128 0 3 0 0 0 4 8 0 0 0 0 0 0 0 86 105 115 105 98 108 101 0 1 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 163 0 0 0 168 0 0 0 4 0 0 2 9 0 0 0 4 0 0 0 9 64 64 128 4 0 128 0 9 64 64 128 4 0 0 1 9 64 64 128 4 0 128 1 9 128 64 128 30 0 128 0 3 0 0 0 4 8 0 0 0 0 0 0 0 86 105 115 105 98 108 101 0 1 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 173 0 0 0 175 0 0 0 2 0 0 6 18 0 0 0 4 0 0 0 69 64 0 0 70 128 192 0 133 192 0 0 196 0 128 0 198 0 193 1 156 128 0 1 197 192 0 0 4 1 128 0 6 1 65 2 220 128 0 1 5 193 0 0 68 1 128 0 70 1 193 2 28 1 0 1 92 128 0 0 9 64 0 128 30 0 128 0 5 0 0 0 4 8 0 0 0 0 0 0 0 65 109 98 105 101 110 116 0 4 7 0 0 0 0 0 0 0 67 111 108 111 114 51 0 4 8 0 0 0 0 0 0 0 102 114 111 109 82 71 66 0 4 9 0 0 0 0 0 0 0 116 111 110 117 109 98 101 114 0 4 5 0 0 0 0 0 0 0 84 101 120 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 205 0 0 0 218 0 0 0 2 4 0 9 32 0 0 0 5 1 0 0 6 65 64 2 65 129 0 0 28 129 0 1 69 1 1 0 70 65 193 2 132 1 0 0 196 1 0 0 4 2 0 0 92 129 0 2 9 65 129 129 9 193 65 131 69 1 1 0 70 65 193 2 128 1 0 0 192 1 128 0 0 2 0 1 92 129 0 2 9 65 1 132 68 1 128 0 9 65 129 132 9 193 0 133 69 193 2 0 70 1 195 2 129 65 3 0 193 65 3 0 1 130 3 0 92 129 0 2 23 64 129 1 22 192 255 127 30 1 0 1 30 0 128 0 15 0 0 0 4 5 0 0 0 0 0 0 0 76 105 109 101 0 4 9 0 0 0 0 0 0 0 67 114 101 97 116 101 85 73 0 4 5 0 0 0 0 0 0 0 80 97 114 116 0 4 5 0 0 0 0 0 0 0 83 105 122 101 0 4 8 0 0 0 0 0 0 0 86 101 99 116 111 114 51 0 4 4 0 0 0 0 0 0 0 110 101 119 0 4 9 0 0 0 0 0 0 0 65 110 99 104 111 114 101 100 0 1 1 4 9 0 0 0 0 0 0 0 80 111 115 105 116 105 111 110 0 4 7 0 0 0 0 0 0 0 80 97 114 101 110 116 0 4 6 0 0 0 0 0 0 0 67 111 108 111 114 0 4 7 0 0 0 0 0 0 0 67 111 108 111 114 51 0 4 8 0 0 0 0 0 0 0 102 114 111 109 82 71 66 0 3 0 0 0 0 0 0 0 0 3 0 0 0 0 0 192 98 64 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 220 0 0 0 242 0 0 0 4 3 0 15 106 0 0 0 197 0 0 0 198 64 192 1 1 129 0 0 65 193 0 0 129 1 1 0 220 128 0 2 5 65 1 0 6 129 65 2 64 1 0 1 28 129 0 1 68 1 0 0 14 65 1 2 68 1 128 0 12 65 1 2 68 1 0 1 24 64 1 2 22 128 1 128 5 1 0 0 6 65 64 2 65 129 0 0 129 129 0 0 193 193 1 0 28 129 0 2 192 0 0 2 4 1 128 1 68 1 0 0 78 65 1 0 133 65 1 0 134 129 65 3 192 1 0 1 156 129 0 1 196 1 0 0 142 193 1 3 196 1 128 0 140 193 1 3 196 1 0 0 206 193 129 0 0 2 128 1 28 129 128 2 68 1 128 0 133 65 1 0 134 129 65 3 192 1 0 1 156 129 0 1 196 1 0 0 142 193 1 3 76 129 129 2 132 1 0 0 77 129 129 2 133 65 1 0 134 129 65 3 192 1 0 1 156 129 0 1 196 1 0 0 142 193 1 3 196 1 128 0 140 193 1 3 196 1 0 1 24 192 1 3 22 128 6 128 132 1 0 1 197 65 1 0 198 129 193 3 0 2 0 1 220 129 0 1 4 2 0 0 206 1 130 3 4 2 128 0 204 1 130 3 24 128 129 3 22 192 3 128 196 1 128 1 4 2 0 0 14 2 2 0 64 2 0 3 132 2 0 0 142 130 130 0 197 2 0 0 198 66 192 5 1 131 0 0 65 131 0 0 129 195 1 0 220 2 0 2 220 65 0 0 196 1 0 0 141 193 1 3 22 64 249 127 24 64 1 129 22 192 3 128 132 1 128 1 196 1 0 0 206 193 1 0 0 2 128 2 68 2 0 0 78 66 130 0 133 2 0 0 134 66 64 5 193 2 2 0 1 3 2 0 65 3 2 0 156 2 0 2 156 65 0 0 132 1 0 0 77 129 129 2 22 64 251 127 30 0 128 0 9 0 0 0 4 7 0 0 0 0 0 0 0 67 111 108 111 114 51 0 4 8 0 0 0 0 0 0 0 102 114 111 109 82 71 66 0 3 0 0 0 0 0 0 0 0 3 0 0 0 0 0 64 99 64 3 0 0 0 0 0 0 55 64 4 5 0 0 0 0 0 0 0 109 97 116 104 0 4 6 0 0 0 0 0 0 0 102 108 111 111 114 0 3 0 0 0 0 0 192 98 64 3 0 0 0 0 0 0 62 64 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 246 0 0 0 5 1 0 0 5 0 0 14 59 0 0 0 5 0 0 0 6 64 64 0 69 128 0 0 90 64 0 0 22 64 0 128 69 192 0 0 92 128 128 0 28 64 0 1 5 0 0 0 6 0 65 0 28 128 128 0 69 0 0 0 70 64 192 0 133 192 0 0 156 0 128 0 92 64 0 0 65 64 1 0 132 0 0 0 193 64 1 0 96 0 9 128 65 65 1 0 132 1 128 0 193 65 1 0 96 1 4 128 69 2 0 0 70 130 193 4 132 2 128 0 143 130 2 4 142 2 0 5 196 2 0 0 207 194 2 2 206 2 128 5 1 195 1 0 92 130 0 2 132 2 0 1 78 130 130 4 132 2 128 1 192 2 0 4 0 3 0 2 64 3 128 4 156 66 0 2 95 65 251 127 68 1 0 2 133 65 2 0 197 1 0 0 198 129 194 3 4 2 0 0 15 2 2 2 14 194 66 4 220 1 0 1 156 129 0 0 193 1 3 0 149 193 1 3 73 129 1 132 69 65 3 0 70 129 195 2 92 65 128 0 95 64 246 127 30 0 128 0 15 0 0 0 4 5 0 0 0 0 0 0 0 109 97 116 104 0 4 11 0 0 0 0 0 0 0 114 97 110 100 111 109 115 101 101 100 0 4 5 0 0 0 0 0 0 0 115 101 101 100 0 4 5 0 0 0 0 0 0 0 116 105 99 107 0 4 7 0 0 0 0 0 0 0 114 97 110 100 111 109 0 3 0 0 0 0 0 0 240 63 4 6 0 0 0 0 0 0 0 110 111 105 115 101 0 3 0 0 0 0 0 0 0 0 4 5 0 0 0 0 0 0 0 84 101 120 116 0 4 9 0 0 0 0 0 0 0 116 111 115 116 114 105 110 103 0 4 6 0 0 0 0 0 0 0 102 108 111 111 114 0 3 0 0 0 0 0 0 89 64 4 2 0 0 0 0 0 0 0 37 0 4 5 0 0 0 0 0 0 0 116 97 115 107 0 4 5 0 0 0 0 0 0 0 119 97 105 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 20 1 0 0 30 1 0 0 5 0 0 7 47 0 0 0 4 0 0 0 11 0 64 0 28 128 0 1 68 0 128 0 134 64 64 0 196 0 0 1 142 192 0 1 76 128 128 0 72 0 128 0 68 0 128 1 134 128 64 0 196 0 0 1 142 192 0 1 76 128 128 0 72 0 128 1 68 0 128 0 24 64 128 129 22 64 0 128 65 192 0 0 72 0 128 0 68 0 128 0 24 0 193 0 22 64 0 128 65 0 1 0 72 0 128 0 68 0 0 2 133 64 1 0 134 128 65 1 196 0 0 2 198 64 193 1 198 192 193 1 156 128 0 1 197 64 1 0 198 0 194 1 5 65 2 0 6 129 66 2 68 1 128 0 28 129 0 1 69 65 2 0 70 129 194 2 132 1 128 1 92 129 0 1 129 193 2 0 220 128 0 2 142 192 0 1 73 128 128 130 30 0 128 0 12 0 0 0 4 14 0 0 0 0 0 0 0 71 101 116 77 111 117 115 101 68 101 108 116 97 0 4 2 0 0 0 0 0 0 0 89 0 4 2 0 0 0 0 0 0 0 88 0 3 0 0 0 0 0 128 86 64 3 0 0 0 0 0 128 86 192 4 7 0 0 0 0 0 0 0 67 70 114 97 109 101 0 4 4 0 0 0 0 0 0 0 110 101 119 0 4 9 0 0 0 0 0 0 0 80 111 115 105 116 105 111 110 0 4 16 0 0 0 0 0 0 0 102 114 111 109 79 114 105 101 110 116 97 116 105 111 110 0 4 5 0 0 0 0 0 0 0 109 97 116 104 0 4 4 0 0 0 0 0 0 0 114 97 100 0 3 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 41 1 0 0 48 1 0 0 4 0 0 5 24 0 0 0 4 0 0 0 6 0 64 0 69 64 0 0 70 0 192 0 70 128 192 0 23 64 0 0 22 192 3 128 4 0 128 0 11 192 64 0 132 0 0 1 134 0 65 1 134 64 65 1 196 0 0 1 198 0 193 1 198 128 193 1 4 1 128 1 206 0 129 1 28 128 0 2 26 0 0 0 22 128 0 128 70 192 65 0 75 0 194 0 92 64 0 1 30 0 128 0 9 0 0 0 4 14 0 0 0 0 0 0 0 77 111 117 115 101 66 101 104 97 118 105 111 114 0 4 5 0 0 0 0 0 0 0 69 110 117 109 0 4 20 0 0 0 0 0 0 0 76 111 99 107 67 117 114 114 101 110 116 80 111 115 105 116 105 111 110 0 4 8 0 0 0 0 0 0 0 82 97 121 99 97 115 116 0 4 7 0 0 0 0 0 0 0 67 70 114 97 109 101 0 4 9 0 0 0 0 0 0 0 80 111 115 105 116 105 111 110 0 4 11 0 0 0 0 0 0 0 76 111 111 107 86 101 99 116 111 114 0 4 9 0 0 0 0 0 0 0 73 110 115 116 97 110 99 101 0 4 8 0 0 0 0 0 0 0 68 101 115 116 114 111 121 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 49 1 0 0 56 1 0 0 5 0 0 11 43 0 0 0 4 0 0 0 11 0 64 0 132 0 128 0 134 64 64 1 134 128 64 1 196 0 128 0 198 64 192 1 198 192 192 1 4 1 0 1 206 0 129 1 28 128 0 2 26 0 0 0 22 0 7 128 69 0 1 0 70 64 193 0 134 128 65 0 134 192 65 1 196 0 128 1 142 192 0 1 198 128 65 0 198 0 194 1 4 1 128 1 206 0 129 1 6 129 65 0 6 65 66 2 68 1 128 1 14 65 1 2 92 128 0 2 134 128 66 0 134 128 64 1 140 64 0 1 196 0 0 2 6 193 65 1 70 1 66 1 134 65 66 1 197 193 2 0 198 1 195 3 1 66 3 0 65 130 3 0 129 194 3 0 220 1 0 2 220 64 0 0 30 0 128 0 16 0 0 0 4 8 0 0 0 0 0 0 0 82 97 121 99 97 115 116 0 4 7 0 0 0 0 0 0 0 67 70 114 97 109 101 0 4 9 0 0 0 0 0 0 0 80 111 115 105 116 105 111 110 0 4 11 0 0 0 0 0 0 0 76 111 111 107 86 101 99 116 111 114 0 4 8 0 0 0 0 0 0 0 86 101 99 116 111 114 51 0 4 4 0 0 0 0 0 0 0 110 101 119 0 4 7 0 0 0 0 0 0 0 78 111 114 109 97 108 0 4 2 0 0 0 0 0 0 0 88 0 4 2 0 0 0 0 0 0 0 89 0 4 2 0 0 0 0 0 0 0 90 0 4 9 0 0 0 0 0 0 0 73 110 115 116 97 110 99 101 0 4 7 0 0 0 0 0 0 0 67 111 108 111 114 51 0 4 8 0 0 0 0 0 0 0 102 114 111 109 82 71 66 0 3 0 0 0 0 0 128 100 64 3 0 0 0 0 0 0 93 64 3 0 0 0 0 0 64 82 64 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 61 1 0 0 75 1 0 0 4 1 0 3 41 0 0 0 70 0 64 0 133 64 0 0 134 0 64 1 134 128 64 1 23 128 128 0 22 64 8 128 68 0 0 0 70 192 192 0 23 0 193 0 22 64 7 128 68 0 128 0 70 64 193 0 133 64 0 0 134 64 65 1 134 128 65 1 23 128 128 0 22 192 2 128 68 0 128 0 133 64 0 0 134 64 65 1 134 192 65 1 73 128 128 130 68 0 128 0 73 64 66 132 68 0 0 1 73 64 194 129 68 0 128 1 73 0 193 129 22 128 2 128 68 0 128 0 133 64 0 0 134 64 65 1 134 128 65 1 73 128 128 130 68 0 128 0 73 0 65 132 68 0 128 1 73 64 194 129 68 0 0 1 73 0 193 129 30 0 128 0 10 0 0 0 4 8 0 0 0 0 0 0 0 75 101 121 67 111 100 101 0 4 5 0 0 0 0 0 0 0 69 110 117 109 0 4 4 0 0 0 0 0 0 0 84 97 98 0 4 8 0 0 0 0 0 0 0 86 105 115 105 98 108 101 0 1 1 4 14 0 0 0 0 0 0 0 77 111 117 115 101 66 101 104 97 118 105 111 114 0 4 8 0 0 0 0 0 0 0 68 101 102 97 117 108 116 0 4 20 0 0 0 0 0 0 0 76 111 99 107 67 117 114 114 101 110 116 80 111 115 105 116 105 111 110 0 4 17 0 0 0 0 0 0 0 77 111 117 115 101 73 99 111 110 69 110 97 98 108 101 100 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 77 1 0 0 83 1 0 0 3 0 0 2 12 0 0 0 4 0 0 0 69 64 0 0 70 0 192 0 70 128 192 0 9 64 0 128 4 0 0 0 9 0 193 129 4 0 128 0 9 128 193 130 4 0 0 1 9 0 193 130 30 0 128 0 7 0 0 0 4 14 0 0 0 0 0 0 0 77 111 117 115 101 66 101 104 97 118 105 111 114 0 4 5 0 0 0 0 0 0 0 69 110 117 109 0 4 20 0 0 0 0 0 0 0 76 111 99 107 67 117 114 114 101 110 116 80 111 115 105 116 105 111 110 0 4 17 0 0 0 0 0 0 0 77 111 117 115 101 73 99 111 110 69 110 97 98 108 101 100 0 1 0 4 8 0 0 0 0 0 0 0 86 105 115 105 98 108 101 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 85 1 0 0 92 1 0 0 6 0 0 3 19 0 0 0 4 0 0 0 11 0 64 0 28 64 0 1 5 64 0 0 6 128 64 0 65 192 0 0 132 0 128 0 28 128 128 1 8 0 0 0 4 0 0 1 11 0 65 0 28 64 0 1 4 0 128 1 9 128 193 130 4 0 0 2 9 128 193 130 4 0 128 2 9 192 193 130 30 0 128 0 8 0 0 0 4 8 0 0 0 0 0 0 0 68 101 115 116 114 111 121 0 4 5 0 0 0 0 0 0 0 76 105 109 101 0 4 9 0 0 0 0 0 0 0 67 114 101 97 116 101 85 73 0 4 7 0 0 0 0 0 0 0 70 111 108 100 101 114 0 4 11 0 0 0 0 0 0 0 68 105 115 99 111 110 110 101 99 116 0 4 8 0 0 0 0 0 0 0 86 105 115 105 98 108 101 0 1 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 98 1 0 0 109 1 0 0 4 1 0 8 45 0 0 0 68 0 0 0 132 0 0 0 134 0 64 1 140 0 0 1 73 128 0 128 68 0 128 0 79 64 192 0 132 0 0 1 77 128 128 0 132 0 128 1 139 128 64 1 5 193 0 0 6 1 65 2 68 1 0 0 70 1 192 2 70 65 193 2 70 129 193 2 132 1 0 0 134 1 64 3 134 65 65 3 134 193 65 3 141 65 0 3 196 1 0 0 198 1 192 3 198 65 193 3 198 1 194 3 28 129 0 2 64 1 0 0 156 128 0 2 154 0 0 0 22 192 2 128 196 0 0 0 4 1 0 0 6 1 64 2 13 1 0 2 201 0 1 128 197 192 0 0 198 0 193 1 1 65 2 0 65 65 2 0 129 65 2 0 221 0 0 2 222 0 0 0 30 0 0 1 30 0 128 0 10 0 0 0 4 7 0 0 0 0 0 0 0 67 70 114 97 109 101 0 3 0 0 0 0 0 0 0 64 4 8 0 0 0 0 0 0 0 82 97 121 99 97 115 116 0 4 8 0 0 0 0 0 0 0 86 101 99 116 111 114 51 0 4 4 0 0 0 0 0 0 0 110 101 119 0 4 9 0 0 0 0 0 0 0 80 111 115 105 116 105 111 110 0 4 2 0 0 0 0 0 0 0 88 0 4 2 0 0 0 0 0 0 0 89 0 4 2 0 0 0 0 0 0 0 90 0 3 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 116 1 0 0 174 1 0 0 13 0 0 4 22 0 0 0 5 0 0 0 6 64 64 0 65 128 0 0 28 128 0 1 70 192 64 0 75 0 193 0 228 0 0 0 4 0 128 0 4 0 0 1 4 0 128 1 4 0 0 2 4 0 128 2 4 0 0 3 4 0 128 3 4 0 0 4 4 0 128 4 4 0 0 5 4 0 128 5 4 0 0 6 92 128 128 1 72 0 0 0 30 0 128 0 5 0 0 0 4 5 0 0 0 0 0 0 0 76 105 109 101 0 4 11 0 0 0 0 0 0 0 71 101 116 83 101 114 118 105 99 101 0 4 11 0 0 0 0 0 0 0 82 117 110 83 101 114 118 105 99 101 0 4 14 0 0 0 0 0 0 0 82 101 110 100 101 114 83 116 101 112 112 101 100 0 4 8 0 0 0 0 0 0 0 67 111 110 110 101 99 116 0 1 0 0 0 0 0 0 0 0 0 0 0 118 1 0 0 173 1 0 0 12 1 0 9 242 0 0 0 68 0 0 0 70 0 192 0 133 64 0 0 134 0 64 1 134 128 64 1 23 128 128 0 22 0 0 128 30 0 128 0 68 0 0 0 75 192 192 0 197 64 0 0 198 0 193 1 198 64 193 1 92 128 128 1 90 0 0 0 22 0 5 128 68 0 128 0 132 0 128 0 134 128 65 1 196 0 0 1 5 193 1 0 6 1 66 2 68 1 128 0 70 129 193 2 70 65 194 2 70 129 194 2 129 193 2 0 196 1 128 0 198 129 193 3 198 65 194 3 198 1 195 3 28 129 0 2 68 1 128 1 14 65 1 2 220 128 0 1 140 192 0 1 73 128 0 131 68 0 0 0 75 192 192 0 197 64 0 0 198 0 193 1 198 64 195 1 92 128 128 1 90 0 0 0 22 64 5 128 68 0 128 0 132 0 128 0 134 128 65 1 196 0 0 1 5 193 1 0 6 1 66 2 68 1 128 0 70 129 193 2 70 65 194 2 70 129 194 2 129 193 2 0 196 1 128 0 198 129 193 3 198 65 194 3 198 1 195 3 28 129 0 2 68 1 128 1 82 1 128 2 14 65 1 2 220 128 0 1 140 192 0 1 73 128 0 131 68 0 0 0 75 192 192 0 197 64 0 0 198 0 193 1 198 128 195 1 92 128 128 1 90 0 0 0 22 192 6 128 68 0 128 0 70 128 193 0 133 128 1 0 134 192 67 1 193 192 2 0 5 1 4 0 6 65 68 2 65 129 4 0 28 129 0 1 65 193 2 0 156 128 0 2 78 128 128 0 70 64 194 0 132 0 128 0 196 0 128 0 198 128 193 1 4 1 0 1 69 193 1 0 70 1 194 2 134 129 194 0 193 193 2 0 6 2 195 0 92 129 0 2 132 1 128 1 78 129 129 2 28 129 0 1 204 0 129 1 137 192 0 131 68 0 0 0 75 192 192 0 197 64 0 0 198 0 193 1 198 192 196 1 92 128 128 1 90 0 0 0 22 192 6 128 68 0 128 0 70 128 193 0 133 128 1 0 134 192 67 1 193 192 2 0 5 1 4 0 6 65 68 2 65 1 5 0 28 129 0 1 65 193 2 0 156 128 0 2 78 128 128 0 70 64 194 0 132 0 128 0 196 0 128 0 198 128 193 1 4 1 0 1 69 193 1 0 70 1 194 2 134 129 194 0 193 193 2 0 6 2 195 0 92 129 0 2 132 1 128 1 78 129 129 2 28 129 0 1 204 0 129 1 137 192 0 131 68 0 0 2 75 64 197 0 196 0 128 0 198 128 193 1 198 128 197 1 5 193 1 0 6 1 66 2 65 193 2 0 132 1 128 2 142 193 69 3 196 1 0 3 140 193 1 3 146 1 0 3 193 193 2 0 28 1 0 2 92 128 0 0 90 64 0 0 22 192 1 128 132 0 128 3 23 192 66 1 22 64 0 128 129 0 6 0 136 0 128 3 130 0 0 0 136 0 0 4 22 64 5 128 130 0 128 0 136 0 0 4 129 192 2 0 136 0 128 3 132 0 128 0 196 0 128 0 198 128 193 1 6 129 197 0 69 193 1 0 70 1 194 2 129 193 2 0 196 1 128 2 206 193 197 3 1 194 2 0 92 129 0 2 12 65 1 2 68 1 128 0 70 129 193 2 70 129 197 2 13 65 1 2 204 0 129 1 137 192 0 131 132 0 0 0 139 192 64 1 5 65 0 0 6 1 65 2 6 65 70 2 156 128 128 1 154 0 0 0 22 0 1 128 132 0 0 4 154 0 0 0 22 64 0 128 129 128 6 0 136 0 128 3 132 0 128 3 87 192 66 1 22 128 6 128 132 0 128 3 24 192 70 1 22 64 0 128 129 192 2 0 136 0 128 3 132 0 128 3 25 192 66 1 22 192 0 128 132 0 128 3 196 0 128 4 140 192 0 1 136 0 128 3 132 0 128 3 196 0 0 5 142 192 0 1 136 0 128 3 132 0 128 0 196 0 128 0 198 128 193 1 5 193 1 0 6 1 66 2 65 193 2 0 132 1 128 3 193 193 2 0 28 129 0 2 204 0 129 1 137 192 0 131 132 0 128 5 197 0 4 0 198 64 199 1 15 1 0 141 220 128 0 1 1 129 7 0 213 0 129 1 137 192 0 142 133 192 7 0 134 0 72 1 156 64 128 0 30 0 128 0 33 0 0 0 4 14 0 0 0 0 0 0 0 77 111 117 115 101 66 101 104 97 118 105 111 114 0 4 5 0 0 0 0 0 0 0 69 110 117 109 0 4 8 0 0 0 0 0 0 0 68 101 102 97 117 108 116 0 4 10 0 0 0 0 0 0 0 73 115 75 101 121 68 111 119 110 0 4 8 0 0 0 0 0 0 0 75 101 121 67 111 100 101 0 4 2 0 0 0 0 0 0 0 87 0 4 7 0 0 0 0 0 0 0 67 70 114 97 109 101 0 4 8 0 0 0 0 0 0 0 86 101 99 116 111 114 51 0 4 4 0 0 0 0 0 0 0 110 101 119 0 4 11 0 0 0 0 0 0 0 76 111 111 107 86 101 99 116 111 114 0 4 2 0 0 0 0 0 0 0 88 0 3 0 0 0 0 0 0 0 0 4 2 0 0 0 0 0 0 0 90 0 4 2 0 0 0 0 0 0 0 83 0 4 2 0 0 0 0 0 0 0 65 0 4 7 0 0 0 0 0 0 0 65 110 103 108 101 115 0 4 5 0 0 0 0 0 0 0 109 97 116 104 0 4 4 0 0 0 0 0 0 0 114 97 100 0 3 0 0 0 0 0 128 86 64 4 2 0 0 0 0 0 0 0 68 0 3 0 0 0 0 0 128 86 192 4 8 0 0 0 0 0 0 0 82 97 121 99 97 115 116 0 4 9 0 0 0 0 0 0 0 80 111 115 105 116 105 111 110 0 3 0 0 0 0 0 0 0 64 3 154 153 153 153 153 153 185 191 4 6 0 0 0 0 0 0 0 83 112 97 99 101 0 3 0 0 0 0 0 0 240 63 3 154 153 153 153 153 153 185 63 4 5 0 0 0 0 0 0 0 84 101 120 116 0 4 6 0 0 0 0 0 0 0 102 108 111 111 114 0 4 5 0 0 0 0 0 0 0 32 70 80 83 0 4 5 0 0 0 0 0 0 0 116 97 115 107 0 4 5 0 0 0 0 0 0 0 119 97 105 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 176 1 0 0 193 1 0 0 8 0 0 6 47 0 0 0 4 0 0 0 9 64 64 128 4 0 128 0 9 64 64 128 4 0 0 1 9 128 64 128 4 0 128 1 9 64 64 128 4 0 0 2 28 64 128 0 5 192 0 0 65 0 1 0 28 64 0 1 4 0 128 2 69 64 1 0 70 128 193 0 133 192 1 0 134 128 65 1 193 0 2 0 1 65 2 0 65 1 2 0 156 0 0 2 92 128 0 0 9 64 128 130 4 0 0 3 69 192 2 0 70 128 194 0 70 0 195 0 9 64 0 133 4 0 0 3 9 64 192 134 5 192 0 0 65 128 3 0 28 64 0 1 4 0 128 3 28 64 128 0 5 192 0 0 65 192 3 0 28 64 0 1 4 0 128 0 9 128 64 128 4 0 0 1 9 64 64 128 5 192 0 0 65 0 4 0 28 64 0 1 30 0 128 0 17 0 0 0 4 8 0 0 0 0 0 0 0 86 105 115 105 98 108 101 0 1 0 1 1 4 4 0 0 0 0 0 0 0 108 111 103 0 4 18 0 0 0 0 0 0 0 116 101 114 114 97 105 110 32 103 101 110 101 114 97 116 101 100 0 4 7 0 0 0 0 0 0 0 67 70 114 97 109 101 0 4 4 0 0 0 0 0 0 0 110 101 119 0 4 8 0 0 0 0 0 0 0 86 101 99 116 111 114 51 0 3 0 0 0 0 0 0 16 64 3 0 0 0 0 0 64 80 64 4 14 0 0 0 0 0 0 0 77 111 117 115 101 66 101 104 97 118 105 111 114 0 4 5 0 0 0 0 0 0 0 69 110 117 109 0 4 20 0 0 0 0 0 0 0 76 111 99 107 67 117 114 114 101 110 116 80 111 115 105 116 105 111 110 0 4 17 0 0 0 0 0 0 0 77 111 117 115 101 73 99 111 110 69 110 97 98 108 101 100 0 4 12 0 0 0 0 0 0 0 99 111 110 102 105 103 32 100 111 110 101 0 4 13 0 0 0 0 0 0 0 114 101 110 100 101 114 32 115 101 116 117 112 0 4 13 0 0 0 0 0 0 0 103 97 109 101 32 118 105 115 105 98 108 101 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 195 1 0 0 201 1 0 0 2 0 0 2 13 0 0 0 5 0 0 0 65 64 0 0 28 64 0 1 4 0 0 0 26 0 0 0 22 128 0 128 4 0 0 0 11 128 64 0 28 64 0 1 4 0 128 0 11 128 64 0 28 64 0 1 30 0 128 0 3 0 0 0 4 4 0 0 0 0 0 0 0 108 111 103 0 4 23 0 0 0 0 0 0 0 98 117 105 108 100 98 114 101 97 107 32 100 105 115 99 111 110 110 101 99 116 115 0 4 11 0 0 0 0 0 0 0 68 105 115 99 111 110 110 101 99 116 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 