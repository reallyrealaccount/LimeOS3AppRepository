LEF            ruben070hallo                   69cc34544e7e8a9a9a9e46322cf95fd3f3bd12104d7b39c8f8c78e9f4cc58423LuaQ         @                @@ A�  ��  ��E   F � �   �@ \���� � B�@ � AA �A ���I� ��� � C�@ A AA �A ���I����� � C�  A A� �� I� ��   � A�   � ����� � �A AA �A �A ܀������� � �� AA �� �A ܀��� ��� � � AA �� ܀ �� ��@E��� ƀ�� ��� ���ƌ� Ǎ��ǎ�� � � AA �� ܀ �����   � �   A� ܀��@I�� CA� �� �� � ��� ��@B���J�    �A�A�J�A    �A���J��  A�  A@  �� ��	�J�E� F��� �� � A� \��	A�E� F��� �A B AB \��	A��	AB�F�IK���     \A�FAJK��    \A�E  F��  �� \���� �C�A B AB �B ���I���IAB�����J$B   ��A��A��J$�   ��A��  �A�  � ����K��� ��� A� �� �� ܁������ ��B AB �B �B ܁������AB���I��d�    �A��AJ��d    �A��  ��   A� ܁��AK�� CA� �� �� � ����� CA� �B �B C ������AB���J�B   �B�B�J��   �B�  A@  �� ��E� F��� �B C AC \��	B��E� F��B �B � AC \��	B�E� F�� �B � \� 	B�	BC�E� F��F�	B�	�ˌ	BB�	B̎	�̍	B̙E� F�� �B � \� 	B�� � 4          Lime        CreateWindow        PhotoLime v1        rbxassetid://9397029482 	       CreateUI        Frame        Size        UDim2 
       fromScale       �?�������?	       Position        new                BackgroundColor3        Color3 �Q���?{�G�z�?       TextButton �������?       BorderSizePixel ������@       Font        Enum        Ubuntu 	       TextSize       D@       Text        Page 1        TextScaled        TextColor3 333333�?�������?      �?       ImageButton        Image +       http://www.roblox.com/asset/?id=8425069718        ZIndex        MouseEnter        Connect        MouseLeave        MouseButton1Click +       http://www.roblox.com/asset/?id=8345858114 +       http://www.roblox.com/asset/?id=8450601351 +       http://www.roblox.com/asset/?id=6075395846 333333�?      6@       BackgroundTransparency         More Soon!        Active                          E@  F�� ��  ��  �  A�  \��	@ �   	@A� �           Size        UDim2        new ��Q��?       ZIndex        @                                                         Image1            "           E@  F�� ��  ��  �  A�  \��	@ �   	@A� �           Size        UDim2        new �������?       ZIndex       �?                                           !   !   "                 Image1         $   &          �            &                   .   1           E@  F�� ��  ��  �  A�  \��	@ �   	@A� �           Size        UDim2        new ��Q��?       ZIndex        @       /   /   /   /   /   /   /   /   /   0   0   1                 Image2         3   6           E@  F�� ��  ��  �  A�  \��	@ �   	@A� �           Size        UDim2        new �������?       ZIndex       �?       4   4   4   4   4   4   4   4   4   5   5   6                 Image2         =   @           E@  F�� ��  ��  �  A�  \��	@ �   	@A� �           Size        UDim2        new ��Q��?       ZIndex        @       >   >   >   >   >   >   >   >   >   ?   ?   @                 Image3         B   E           E@  F�� ��  ��  �  A�  \��	@ �   	@A� �           Size        UDim2        new �������?       ZIndex       �?       C   C   C   C   C   C   C   C   C   D   D   E                 Image3         N   Q           E@  F�� ��  ��  �  A�  \��	@ �   	@A� �           Size        UDim2        new ��Q��?       ZIndex        @       O   O   O   O   O   O   O   O   O   P   P   Q                 Image4         S   V           E@  F�� ��  ��  �  A�  \��	@ �   	@A� �           Size        UDim2        new �������?       ZIndex       �?       T   T   T   T   T   T   T   T   T   U   U   V                 Image4         _   b           E@  F�� ��  ��  �  A�  \��	@ �   	@A� �           Size        UDim2        new ��Q��?       ZIndex        @       `   `   `   `   `   `   `   `   `   a   a   b                 Image5         d   g           E@  F�� ��  ��  �  A�  \��	@ �   	@A� �           Size        UDim2        new �������?       ZIndex       �?       e   e   e   e   e   e   e   e   e   f   f   g                 Image5                                                                                                      
   
   
   
   
                                                                                                                                                                                       "   "      $   $   &   $   (   (   (   (   (   )   *   *   *   *   *   *   *   *   +   +   +   +   +   +   +   +   ,   .   .   1   1   .   3   3   6   6   3   8   8   8   8   8   :   :   :   :   :   :   :   :   ;   =   =   @   @   =   B   B   E   E   B   H   H   H   H   H   I   J   J   J   J   J   J   J   J   K   K   K   K   K   K   K   K   L   N   N   Q   Q   N   S   S   V   V   S   Y   Y   Y   Y   Y   Z   [   [   [   [   [   [   [   [   \   \   \   \   \   \   \   \   ]   _   _   b   b   _   d   d   g   g   d   i   i   i   i   i   j   j   j   j   j   j   j   j   k   k   k   k   k   k   k   k   l   l   l   l   l   l   l   m   n   n   n   n   o   p   q   r   s   u   u   u   u   u   u   u   u   	          app             bar 
            HomeButton &            Image1 Q            Image2 n            Image3 �            Image4 �            Image5 �            HomeButton2 �         